magic
tech sky130A
magscale 1 2
timestamp 1654747626
<< obsli1 >>
rect 1104 2159 213532 214353
<< obsm1 >>
rect 566 484 214438 214464
<< metal2 >>
rect 938 215988 994 216788
rect 2778 215988 2834 216788
rect 4618 215988 4674 216788
rect 6550 215988 6606 216788
rect 8390 215988 8446 216788
rect 10322 215988 10378 216788
rect 12162 215988 12218 216788
rect 14094 215988 14150 216788
rect 15934 215988 15990 216788
rect 17866 215988 17922 216788
rect 19706 215988 19762 216788
rect 21638 215988 21694 216788
rect 23478 215988 23534 216788
rect 25410 215988 25466 216788
rect 27250 215988 27306 216788
rect 29090 215988 29146 216788
rect 31022 215988 31078 216788
rect 32862 215988 32918 216788
rect 34794 215988 34850 216788
rect 36634 215988 36690 216788
rect 38566 215988 38622 216788
rect 40406 215988 40462 216788
rect 42338 215988 42394 216788
rect 44178 215988 44234 216788
rect 46110 215988 46166 216788
rect 47950 215988 48006 216788
rect 49882 215988 49938 216788
rect 51722 215988 51778 216788
rect 53654 215988 53710 216788
rect 55494 215988 55550 216788
rect 57334 215988 57390 216788
rect 59266 215988 59322 216788
rect 61106 215988 61162 216788
rect 63038 215988 63094 216788
rect 64878 215988 64934 216788
rect 66810 215988 66866 216788
rect 68650 215988 68706 216788
rect 70582 215988 70638 216788
rect 72422 215988 72478 216788
rect 74354 215988 74410 216788
rect 76194 215988 76250 216788
rect 78126 215988 78182 216788
rect 79966 215988 80022 216788
rect 81806 215988 81862 216788
rect 83738 215988 83794 216788
rect 85578 215988 85634 216788
rect 87510 215988 87566 216788
rect 89350 215988 89406 216788
rect 91282 215988 91338 216788
rect 93122 215988 93178 216788
rect 95054 215988 95110 216788
rect 96894 215988 96950 216788
rect 98826 215988 98882 216788
rect 100666 215988 100722 216788
rect 102598 215988 102654 216788
rect 104438 215988 104494 216788
rect 106370 215988 106426 216788
rect 108210 215988 108266 216788
rect 110050 215988 110106 216788
rect 111982 215988 112038 216788
rect 113822 215988 113878 216788
rect 115754 215988 115810 216788
rect 117594 215988 117650 216788
rect 119526 215988 119582 216788
rect 121366 215988 121422 216788
rect 123298 215988 123354 216788
rect 125138 215988 125194 216788
rect 127070 215988 127126 216788
rect 128910 215988 128966 216788
rect 130842 215988 130898 216788
rect 132682 215988 132738 216788
rect 134614 215988 134670 216788
rect 136454 215988 136510 216788
rect 138294 215988 138350 216788
rect 140226 215988 140282 216788
rect 142066 215988 142122 216788
rect 143998 215988 144054 216788
rect 145838 215988 145894 216788
rect 147770 215988 147826 216788
rect 149610 215988 149666 216788
rect 151542 215988 151598 216788
rect 153382 215988 153438 216788
rect 155314 215988 155370 216788
rect 157154 215988 157210 216788
rect 159086 215988 159142 216788
rect 160926 215988 160982 216788
rect 162766 215988 162822 216788
rect 164698 215988 164754 216788
rect 166538 215988 166594 216788
rect 168470 215988 168526 216788
rect 170310 215988 170366 216788
rect 172242 215988 172298 216788
rect 174082 215988 174138 216788
rect 176014 215988 176070 216788
rect 177854 215988 177910 216788
rect 179786 215988 179842 216788
rect 181626 215988 181682 216788
rect 183558 215988 183614 216788
rect 185398 215988 185454 216788
rect 187330 215988 187386 216788
rect 189170 215988 189226 216788
rect 191010 215988 191066 216788
rect 192942 215988 192998 216788
rect 194782 215988 194838 216788
rect 196714 215988 196770 216788
rect 198554 215988 198610 216788
rect 200486 215988 200542 216788
rect 202326 215988 202382 216788
rect 204258 215988 204314 216788
rect 206098 215988 206154 216788
rect 208030 215988 208086 216788
rect 209870 215988 209926 216788
rect 211802 215988 211858 216788
rect 213642 215988 213698 216788
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8850 0 8906 800
rect 9310 0 9366 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21914 0 21970 800
rect 22374 0 22430 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25410 0 25466 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30194 0 30250 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31482 0 31538 800
rect 31942 0 31998 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33230 0 33286 800
rect 33690 0 33746 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 38014 0 38070 800
rect 38474 0 38530 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41510 0 41566 800
rect 41970 0 42026 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46294 0 46350 800
rect 46754 0 46810 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 48042 0 48098 800
rect 48502 0 48558 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49790 0 49846 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54574 0 54630 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56322 0 56378 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57610 0 57666 800
rect 58070 0 58126 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61106 0 61162 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62394 0 62450 800
rect 62854 0 62910 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64602 0 64658 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65890 0 65946 800
rect 66350 0 66406 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 68466 0 68522 800
rect 68926 0 68982 800
rect 69386 0 69442 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70674 0 70730 800
rect 71134 0 71190 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72422 0 72478 800
rect 72882 0 72938 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 74170 0 74226 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77206 0 77262 800
rect 77666 0 77722 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78954 0 79010 800
rect 79414 0 79470 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80702 0 80758 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81990 0 82046 800
rect 82450 0 82506 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83738 0 83794 800
rect 84198 0 84254 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85486 0 85542 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86774 0 86830 800
rect 87234 0 87290 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88522 0 88578 800
rect 88982 0 89038 800
rect 89442 0 89498 800
rect 89810 0 89866 800
rect 90270 0 90326 800
rect 90730 0 90786 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93306 0 93362 800
rect 93766 0 93822 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 95054 0 95110 800
rect 95514 0 95570 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96802 0 96858 800
rect 97262 0 97318 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98550 0 98606 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99838 0 99894 800
rect 100298 0 100354 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101586 0 101642 800
rect 102046 0 102102 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103334 0 103390 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 105082 0 105138 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106370 0 106426 800
rect 106830 0 106886 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 108118 0 108174 800
rect 108578 0 108634 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109866 0 109922 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112902 0 112958 800
rect 113362 0 113418 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114650 0 114706 800
rect 115110 0 115166 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117686 0 117742 800
rect 118146 0 118202 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119434 0 119490 800
rect 119894 0 119950 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121182 0 121238 800
rect 121642 0 121698 800
rect 122102 0 122158 800
rect 122470 0 122526 800
rect 122930 0 122986 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124218 0 124274 800
rect 124678 0 124734 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125966 0 126022 800
rect 126426 0 126482 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127714 0 127770 800
rect 128174 0 128230 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129462 0 129518 800
rect 129922 0 129978 800
rect 130290 0 130346 800
rect 130750 0 130806 800
rect 131210 0 131266 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132498 0 132554 800
rect 132958 0 133014 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134246 0 134302 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135534 0 135590 800
rect 135994 0 136050 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137282 0 137338 800
rect 137742 0 137798 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 139030 0 139086 800
rect 139490 0 139546 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140778 0 140834 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 142066 0 142122 800
rect 142526 0 142582 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143814 0 143870 800
rect 144274 0 144330 800
rect 144734 0 144790 800
rect 145102 0 145158 800
rect 145562 0 145618 800
rect 146022 0 146078 800
rect 146482 0 146538 800
rect 146850 0 146906 800
rect 147310 0 147366 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148598 0 148654 800
rect 149058 0 149114 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150346 0 150402 800
rect 150806 0 150862 800
rect 151266 0 151322 800
rect 151634 0 151690 800
rect 152094 0 152150 800
rect 152554 0 152610 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153842 0 153898 800
rect 154302 0 154358 800
rect 154670 0 154726 800
rect 155130 0 155186 800
rect 155590 0 155646 800
rect 156050 0 156106 800
rect 156418 0 156474 800
rect 156878 0 156934 800
rect 157338 0 157394 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158626 0 158682 800
rect 159086 0 159142 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160374 0 160430 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161662 0 161718 800
rect 162122 0 162178 800
rect 162582 0 162638 800
rect 162950 0 163006 800
rect 163410 0 163466 800
rect 163870 0 163926 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165158 0 165214 800
rect 165618 0 165674 800
rect 165986 0 166042 800
rect 166446 0 166502 800
rect 166906 0 166962 800
rect 167366 0 167422 800
rect 167734 0 167790 800
rect 168194 0 168250 800
rect 168654 0 168710 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169942 0 169998 800
rect 170402 0 170458 800
rect 170862 0 170918 800
rect 171230 0 171286 800
rect 171690 0 171746 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172978 0 173034 800
rect 173438 0 173494 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174726 0 174782 800
rect 175186 0 175242 800
rect 175646 0 175702 800
rect 176014 0 176070 800
rect 176474 0 176530 800
rect 176934 0 176990 800
rect 177394 0 177450 800
rect 177762 0 177818 800
rect 178222 0 178278 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179510 0 179566 800
rect 179970 0 180026 800
rect 180430 0 180486 800
rect 180798 0 180854 800
rect 181258 0 181314 800
rect 181718 0 181774 800
rect 182178 0 182234 800
rect 182546 0 182602 800
rect 183006 0 183062 800
rect 183466 0 183522 800
rect 183926 0 183982 800
rect 184294 0 184350 800
rect 184754 0 184810 800
rect 185214 0 185270 800
rect 185582 0 185638 800
rect 186042 0 186098 800
rect 186502 0 186558 800
rect 186962 0 187018 800
rect 187330 0 187386 800
rect 187790 0 187846 800
rect 188250 0 188306 800
rect 188710 0 188766 800
rect 189078 0 189134 800
rect 189538 0 189594 800
rect 189998 0 190054 800
rect 190366 0 190422 800
rect 190826 0 190882 800
rect 191286 0 191342 800
rect 191746 0 191802 800
rect 192114 0 192170 800
rect 192574 0 192630 800
rect 193034 0 193090 800
rect 193494 0 193550 800
rect 193862 0 193918 800
rect 194322 0 194378 800
rect 194782 0 194838 800
rect 195242 0 195298 800
rect 195610 0 195666 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 196898 0 196954 800
rect 197358 0 197414 800
rect 197818 0 197874 800
rect 198278 0 198334 800
rect 198646 0 198702 800
rect 199106 0 199162 800
rect 199566 0 199622 800
rect 200026 0 200082 800
rect 200394 0 200450 800
rect 200854 0 200910 800
rect 201314 0 201370 800
rect 201774 0 201830 800
rect 202142 0 202198 800
rect 202602 0 202658 800
rect 203062 0 203118 800
rect 203430 0 203486 800
rect 203890 0 203946 800
rect 204350 0 204406 800
rect 204810 0 204866 800
rect 205178 0 205234 800
rect 205638 0 205694 800
rect 206098 0 206154 800
rect 206558 0 206614 800
rect 206926 0 206982 800
rect 207386 0 207442 800
rect 207846 0 207902 800
rect 208306 0 208362 800
rect 208674 0 208730 800
rect 209134 0 209190 800
rect 209594 0 209650 800
rect 209962 0 210018 800
rect 210422 0 210478 800
rect 210882 0 210938 800
rect 211342 0 211398 800
rect 211710 0 211766 800
rect 212170 0 212226 800
rect 212630 0 212686 800
rect 213090 0 213146 800
rect 213458 0 213514 800
rect 213918 0 213974 800
rect 214378 0 214434 800
<< obsm2 >>
rect 202 215932 882 216050
rect 1050 215932 2722 216050
rect 2890 215932 4562 216050
rect 4730 215932 6494 216050
rect 6662 215932 8334 216050
rect 8502 215932 10266 216050
rect 10434 215932 12106 216050
rect 12274 215932 14038 216050
rect 14206 215932 15878 216050
rect 16046 215932 17810 216050
rect 17978 215932 19650 216050
rect 19818 215932 21582 216050
rect 21750 215932 23422 216050
rect 23590 215932 25354 216050
rect 25522 215932 27194 216050
rect 27362 215932 29034 216050
rect 29202 215932 30966 216050
rect 31134 215932 32806 216050
rect 32974 215932 34738 216050
rect 34906 215932 36578 216050
rect 36746 215932 38510 216050
rect 38678 215932 40350 216050
rect 40518 215932 42282 216050
rect 42450 215932 44122 216050
rect 44290 215932 46054 216050
rect 46222 215932 47894 216050
rect 48062 215932 49826 216050
rect 49994 215932 51666 216050
rect 51834 215932 53598 216050
rect 53766 215932 55438 216050
rect 55606 215932 57278 216050
rect 57446 215932 59210 216050
rect 59378 215932 61050 216050
rect 61218 215932 62982 216050
rect 63150 215932 64822 216050
rect 64990 215932 66754 216050
rect 66922 215932 68594 216050
rect 68762 215932 70526 216050
rect 70694 215932 72366 216050
rect 72534 215932 74298 216050
rect 74466 215932 76138 216050
rect 76306 215932 78070 216050
rect 78238 215932 79910 216050
rect 80078 215932 81750 216050
rect 81918 215932 83682 216050
rect 83850 215932 85522 216050
rect 85690 215932 87454 216050
rect 87622 215932 89294 216050
rect 89462 215932 91226 216050
rect 91394 215932 93066 216050
rect 93234 215932 94998 216050
rect 95166 215932 96838 216050
rect 97006 215932 98770 216050
rect 98938 215932 100610 216050
rect 100778 215932 102542 216050
rect 102710 215932 104382 216050
rect 104550 215932 106314 216050
rect 106482 215932 108154 216050
rect 108322 215932 109994 216050
rect 110162 215932 111926 216050
rect 112094 215932 113766 216050
rect 113934 215932 115698 216050
rect 115866 215932 117538 216050
rect 117706 215932 119470 216050
rect 119638 215932 121310 216050
rect 121478 215932 123242 216050
rect 123410 215932 125082 216050
rect 125250 215932 127014 216050
rect 127182 215932 128854 216050
rect 129022 215932 130786 216050
rect 130954 215932 132626 216050
rect 132794 215932 134558 216050
rect 134726 215932 136398 216050
rect 136566 215932 138238 216050
rect 138406 215932 140170 216050
rect 140338 215932 142010 216050
rect 142178 215932 143942 216050
rect 144110 215932 145782 216050
rect 145950 215932 147714 216050
rect 147882 215932 149554 216050
rect 149722 215932 151486 216050
rect 151654 215932 153326 216050
rect 153494 215932 155258 216050
rect 155426 215932 157098 216050
rect 157266 215932 159030 216050
rect 159198 215932 160870 216050
rect 161038 215932 162710 216050
rect 162878 215932 164642 216050
rect 164810 215932 166482 216050
rect 166650 215932 168414 216050
rect 168582 215932 170254 216050
rect 170422 215932 172186 216050
rect 172354 215932 174026 216050
rect 174194 215932 175958 216050
rect 176126 215932 177798 216050
rect 177966 215932 179730 216050
rect 179898 215932 181570 216050
rect 181738 215932 183502 216050
rect 183670 215932 185342 216050
rect 185510 215932 187274 216050
rect 187442 215932 189114 216050
rect 189282 215932 190954 216050
rect 191122 215932 192886 216050
rect 193054 215932 194726 216050
rect 194894 215932 196658 216050
rect 196826 215932 198498 216050
rect 198666 215932 200430 216050
rect 200598 215932 202270 216050
rect 202438 215932 204202 216050
rect 204370 215932 206042 216050
rect 206210 215932 207974 216050
rect 208142 215932 209814 216050
rect 209982 215932 211746 216050
rect 211914 215932 213586 216050
rect 213754 215932 214432 216050
rect 202 856 214432 215932
rect 314 478 514 856
rect 682 478 974 856
rect 1142 478 1434 856
rect 1602 478 1802 856
rect 1970 478 2262 856
rect 2430 478 2722 856
rect 2890 478 3182 856
rect 3350 478 3550 856
rect 3718 478 4010 856
rect 4178 478 4470 856
rect 4638 478 4930 856
rect 5098 478 5298 856
rect 5466 478 5758 856
rect 5926 478 6218 856
rect 6386 478 6586 856
rect 6754 478 7046 856
rect 7214 478 7506 856
rect 7674 478 7966 856
rect 8134 478 8334 856
rect 8502 478 8794 856
rect 8962 478 9254 856
rect 9422 478 9714 856
rect 9882 478 10082 856
rect 10250 478 10542 856
rect 10710 478 11002 856
rect 11170 478 11462 856
rect 11630 478 11830 856
rect 11998 478 12290 856
rect 12458 478 12750 856
rect 12918 478 13118 856
rect 13286 478 13578 856
rect 13746 478 14038 856
rect 14206 478 14498 856
rect 14666 478 14866 856
rect 15034 478 15326 856
rect 15494 478 15786 856
rect 15954 478 16246 856
rect 16414 478 16614 856
rect 16782 478 17074 856
rect 17242 478 17534 856
rect 17702 478 17994 856
rect 18162 478 18362 856
rect 18530 478 18822 856
rect 18990 478 19282 856
rect 19450 478 19650 856
rect 19818 478 20110 856
rect 20278 478 20570 856
rect 20738 478 21030 856
rect 21198 478 21398 856
rect 21566 478 21858 856
rect 22026 478 22318 856
rect 22486 478 22778 856
rect 22946 478 23146 856
rect 23314 478 23606 856
rect 23774 478 24066 856
rect 24234 478 24526 856
rect 24694 478 24894 856
rect 25062 478 25354 856
rect 25522 478 25814 856
rect 25982 478 26182 856
rect 26350 478 26642 856
rect 26810 478 27102 856
rect 27270 478 27562 856
rect 27730 478 27930 856
rect 28098 478 28390 856
rect 28558 478 28850 856
rect 29018 478 29310 856
rect 29478 478 29678 856
rect 29846 478 30138 856
rect 30306 478 30598 856
rect 30766 478 30966 856
rect 31134 478 31426 856
rect 31594 478 31886 856
rect 32054 478 32346 856
rect 32514 478 32714 856
rect 32882 478 33174 856
rect 33342 478 33634 856
rect 33802 478 34094 856
rect 34262 478 34462 856
rect 34630 478 34922 856
rect 35090 478 35382 856
rect 35550 478 35842 856
rect 36010 478 36210 856
rect 36378 478 36670 856
rect 36838 478 37130 856
rect 37298 478 37498 856
rect 37666 478 37958 856
rect 38126 478 38418 856
rect 38586 478 38878 856
rect 39046 478 39246 856
rect 39414 478 39706 856
rect 39874 478 40166 856
rect 40334 478 40626 856
rect 40794 478 40994 856
rect 41162 478 41454 856
rect 41622 478 41914 856
rect 42082 478 42374 856
rect 42542 478 42742 856
rect 42910 478 43202 856
rect 43370 478 43662 856
rect 43830 478 44030 856
rect 44198 478 44490 856
rect 44658 478 44950 856
rect 45118 478 45410 856
rect 45578 478 45778 856
rect 45946 478 46238 856
rect 46406 478 46698 856
rect 46866 478 47158 856
rect 47326 478 47526 856
rect 47694 478 47986 856
rect 48154 478 48446 856
rect 48614 478 48906 856
rect 49074 478 49274 856
rect 49442 478 49734 856
rect 49902 478 50194 856
rect 50362 478 50562 856
rect 50730 478 51022 856
rect 51190 478 51482 856
rect 51650 478 51942 856
rect 52110 478 52310 856
rect 52478 478 52770 856
rect 52938 478 53230 856
rect 53398 478 53690 856
rect 53858 478 54058 856
rect 54226 478 54518 856
rect 54686 478 54978 856
rect 55146 478 55346 856
rect 55514 478 55806 856
rect 55974 478 56266 856
rect 56434 478 56726 856
rect 56894 478 57094 856
rect 57262 478 57554 856
rect 57722 478 58014 856
rect 58182 478 58474 856
rect 58642 478 58842 856
rect 59010 478 59302 856
rect 59470 478 59762 856
rect 59930 478 60222 856
rect 60390 478 60590 856
rect 60758 478 61050 856
rect 61218 478 61510 856
rect 61678 478 61878 856
rect 62046 478 62338 856
rect 62506 478 62798 856
rect 62966 478 63258 856
rect 63426 478 63626 856
rect 63794 478 64086 856
rect 64254 478 64546 856
rect 64714 478 65006 856
rect 65174 478 65374 856
rect 65542 478 65834 856
rect 66002 478 66294 856
rect 66462 478 66754 856
rect 66922 478 67122 856
rect 67290 478 67582 856
rect 67750 478 68042 856
rect 68210 478 68410 856
rect 68578 478 68870 856
rect 69038 478 69330 856
rect 69498 478 69790 856
rect 69958 478 70158 856
rect 70326 478 70618 856
rect 70786 478 71078 856
rect 71246 478 71538 856
rect 71706 478 71906 856
rect 72074 478 72366 856
rect 72534 478 72826 856
rect 72994 478 73286 856
rect 73454 478 73654 856
rect 73822 478 74114 856
rect 74282 478 74574 856
rect 74742 478 74942 856
rect 75110 478 75402 856
rect 75570 478 75862 856
rect 76030 478 76322 856
rect 76490 478 76690 856
rect 76858 478 77150 856
rect 77318 478 77610 856
rect 77778 478 78070 856
rect 78238 478 78438 856
rect 78606 478 78898 856
rect 79066 478 79358 856
rect 79526 478 79818 856
rect 79986 478 80186 856
rect 80354 478 80646 856
rect 80814 478 81106 856
rect 81274 478 81474 856
rect 81642 478 81934 856
rect 82102 478 82394 856
rect 82562 478 82854 856
rect 83022 478 83222 856
rect 83390 478 83682 856
rect 83850 478 84142 856
rect 84310 478 84602 856
rect 84770 478 84970 856
rect 85138 478 85430 856
rect 85598 478 85890 856
rect 86058 478 86258 856
rect 86426 478 86718 856
rect 86886 478 87178 856
rect 87346 478 87638 856
rect 87806 478 88006 856
rect 88174 478 88466 856
rect 88634 478 88926 856
rect 89094 478 89386 856
rect 89554 478 89754 856
rect 89922 478 90214 856
rect 90382 478 90674 856
rect 90842 478 91134 856
rect 91302 478 91502 856
rect 91670 478 91962 856
rect 92130 478 92422 856
rect 92590 478 92790 856
rect 92958 478 93250 856
rect 93418 478 93710 856
rect 93878 478 94170 856
rect 94338 478 94538 856
rect 94706 478 94998 856
rect 95166 478 95458 856
rect 95626 478 95918 856
rect 96086 478 96286 856
rect 96454 478 96746 856
rect 96914 478 97206 856
rect 97374 478 97666 856
rect 97834 478 98034 856
rect 98202 478 98494 856
rect 98662 478 98954 856
rect 99122 478 99322 856
rect 99490 478 99782 856
rect 99950 478 100242 856
rect 100410 478 100702 856
rect 100870 478 101070 856
rect 101238 478 101530 856
rect 101698 478 101990 856
rect 102158 478 102450 856
rect 102618 478 102818 856
rect 102986 478 103278 856
rect 103446 478 103738 856
rect 103906 478 104198 856
rect 104366 478 104566 856
rect 104734 478 105026 856
rect 105194 478 105486 856
rect 105654 478 105854 856
rect 106022 478 106314 856
rect 106482 478 106774 856
rect 106942 478 107234 856
rect 107402 478 107602 856
rect 107770 478 108062 856
rect 108230 478 108522 856
rect 108690 478 108982 856
rect 109150 478 109350 856
rect 109518 478 109810 856
rect 109978 478 110270 856
rect 110438 478 110638 856
rect 110806 478 111098 856
rect 111266 478 111558 856
rect 111726 478 112018 856
rect 112186 478 112386 856
rect 112554 478 112846 856
rect 113014 478 113306 856
rect 113474 478 113766 856
rect 113934 478 114134 856
rect 114302 478 114594 856
rect 114762 478 115054 856
rect 115222 478 115514 856
rect 115682 478 115882 856
rect 116050 478 116342 856
rect 116510 478 116802 856
rect 116970 478 117170 856
rect 117338 478 117630 856
rect 117798 478 118090 856
rect 118258 478 118550 856
rect 118718 478 118918 856
rect 119086 478 119378 856
rect 119546 478 119838 856
rect 120006 478 120298 856
rect 120466 478 120666 856
rect 120834 478 121126 856
rect 121294 478 121586 856
rect 121754 478 122046 856
rect 122214 478 122414 856
rect 122582 478 122874 856
rect 123042 478 123334 856
rect 123502 478 123702 856
rect 123870 478 124162 856
rect 124330 478 124622 856
rect 124790 478 125082 856
rect 125250 478 125450 856
rect 125618 478 125910 856
rect 126078 478 126370 856
rect 126538 478 126830 856
rect 126998 478 127198 856
rect 127366 478 127658 856
rect 127826 478 128118 856
rect 128286 478 128578 856
rect 128746 478 128946 856
rect 129114 478 129406 856
rect 129574 478 129866 856
rect 130034 478 130234 856
rect 130402 478 130694 856
rect 130862 478 131154 856
rect 131322 478 131614 856
rect 131782 478 131982 856
rect 132150 478 132442 856
rect 132610 478 132902 856
rect 133070 478 133362 856
rect 133530 478 133730 856
rect 133898 478 134190 856
rect 134358 478 134650 856
rect 134818 478 135018 856
rect 135186 478 135478 856
rect 135646 478 135938 856
rect 136106 478 136398 856
rect 136566 478 136766 856
rect 136934 478 137226 856
rect 137394 478 137686 856
rect 137854 478 138146 856
rect 138314 478 138514 856
rect 138682 478 138974 856
rect 139142 478 139434 856
rect 139602 478 139894 856
rect 140062 478 140262 856
rect 140430 478 140722 856
rect 140890 478 141182 856
rect 141350 478 141550 856
rect 141718 478 142010 856
rect 142178 478 142470 856
rect 142638 478 142930 856
rect 143098 478 143298 856
rect 143466 478 143758 856
rect 143926 478 144218 856
rect 144386 478 144678 856
rect 144846 478 145046 856
rect 145214 478 145506 856
rect 145674 478 145966 856
rect 146134 478 146426 856
rect 146594 478 146794 856
rect 146962 478 147254 856
rect 147422 478 147714 856
rect 147882 478 148082 856
rect 148250 478 148542 856
rect 148710 478 149002 856
rect 149170 478 149462 856
rect 149630 478 149830 856
rect 149998 478 150290 856
rect 150458 478 150750 856
rect 150918 478 151210 856
rect 151378 478 151578 856
rect 151746 478 152038 856
rect 152206 478 152498 856
rect 152666 478 152958 856
rect 153126 478 153326 856
rect 153494 478 153786 856
rect 153954 478 154246 856
rect 154414 478 154614 856
rect 154782 478 155074 856
rect 155242 478 155534 856
rect 155702 478 155994 856
rect 156162 478 156362 856
rect 156530 478 156822 856
rect 156990 478 157282 856
rect 157450 478 157742 856
rect 157910 478 158110 856
rect 158278 478 158570 856
rect 158738 478 159030 856
rect 159198 478 159490 856
rect 159658 478 159858 856
rect 160026 478 160318 856
rect 160486 478 160778 856
rect 160946 478 161146 856
rect 161314 478 161606 856
rect 161774 478 162066 856
rect 162234 478 162526 856
rect 162694 478 162894 856
rect 163062 478 163354 856
rect 163522 478 163814 856
rect 163982 478 164274 856
rect 164442 478 164642 856
rect 164810 478 165102 856
rect 165270 478 165562 856
rect 165730 478 165930 856
rect 166098 478 166390 856
rect 166558 478 166850 856
rect 167018 478 167310 856
rect 167478 478 167678 856
rect 167846 478 168138 856
rect 168306 478 168598 856
rect 168766 478 169058 856
rect 169226 478 169426 856
rect 169594 478 169886 856
rect 170054 478 170346 856
rect 170514 478 170806 856
rect 170974 478 171174 856
rect 171342 478 171634 856
rect 171802 478 172094 856
rect 172262 478 172462 856
rect 172630 478 172922 856
rect 173090 478 173382 856
rect 173550 478 173842 856
rect 174010 478 174210 856
rect 174378 478 174670 856
rect 174838 478 175130 856
rect 175298 478 175590 856
rect 175758 478 175958 856
rect 176126 478 176418 856
rect 176586 478 176878 856
rect 177046 478 177338 856
rect 177506 478 177706 856
rect 177874 478 178166 856
rect 178334 478 178626 856
rect 178794 478 178994 856
rect 179162 478 179454 856
rect 179622 478 179914 856
rect 180082 478 180374 856
rect 180542 478 180742 856
rect 180910 478 181202 856
rect 181370 478 181662 856
rect 181830 478 182122 856
rect 182290 478 182490 856
rect 182658 478 182950 856
rect 183118 478 183410 856
rect 183578 478 183870 856
rect 184038 478 184238 856
rect 184406 478 184698 856
rect 184866 478 185158 856
rect 185326 478 185526 856
rect 185694 478 185986 856
rect 186154 478 186446 856
rect 186614 478 186906 856
rect 187074 478 187274 856
rect 187442 478 187734 856
rect 187902 478 188194 856
rect 188362 478 188654 856
rect 188822 478 189022 856
rect 189190 478 189482 856
rect 189650 478 189942 856
rect 190110 478 190310 856
rect 190478 478 190770 856
rect 190938 478 191230 856
rect 191398 478 191690 856
rect 191858 478 192058 856
rect 192226 478 192518 856
rect 192686 478 192978 856
rect 193146 478 193438 856
rect 193606 478 193806 856
rect 193974 478 194266 856
rect 194434 478 194726 856
rect 194894 478 195186 856
rect 195354 478 195554 856
rect 195722 478 196014 856
rect 196182 478 196474 856
rect 196642 478 196842 856
rect 197010 478 197302 856
rect 197470 478 197762 856
rect 197930 478 198222 856
rect 198390 478 198590 856
rect 198758 478 199050 856
rect 199218 478 199510 856
rect 199678 478 199970 856
rect 200138 478 200338 856
rect 200506 478 200798 856
rect 200966 478 201258 856
rect 201426 478 201718 856
rect 201886 478 202086 856
rect 202254 478 202546 856
rect 202714 478 203006 856
rect 203174 478 203374 856
rect 203542 478 203834 856
rect 204002 478 204294 856
rect 204462 478 204754 856
rect 204922 478 205122 856
rect 205290 478 205582 856
rect 205750 478 206042 856
rect 206210 478 206502 856
rect 206670 478 206870 856
rect 207038 478 207330 856
rect 207498 478 207790 856
rect 207958 478 208250 856
rect 208418 478 208618 856
rect 208786 478 209078 856
rect 209246 478 209538 856
rect 209706 478 209906 856
rect 210074 478 210366 856
rect 210534 478 210826 856
rect 210994 478 211286 856
rect 211454 478 211654 856
rect 211822 478 212114 856
rect 212282 478 212574 856
rect 212742 478 213034 856
rect 213202 478 213402 856
rect 213570 478 213862 856
rect 214030 478 214322 856
<< obsm3 >>
rect 197 851 204208 214369
<< metal4 >>
rect 4208 2128 4528 214384
rect 19568 2128 19888 214384
rect 34928 2128 35248 214384
rect 50288 2128 50608 214384
rect 65648 2128 65968 214384
rect 81008 2128 81328 214384
rect 96368 2128 96688 214384
rect 111728 2128 112048 214384
rect 127088 2128 127408 214384
rect 142448 2128 142768 214384
rect 157808 2128 158128 214384
rect 173168 2128 173488 214384
rect 188528 2128 188848 214384
rect 203888 2128 204208 214384
<< obsm4 >>
rect 19379 2347 19488 214029
rect 19968 2347 34848 214029
rect 35328 2347 50208 214029
rect 50688 2347 65568 214029
rect 66048 2347 80928 214029
rect 81408 2347 96288 214029
rect 96768 2347 111648 214029
rect 112128 2347 127008 214029
rect 127488 2347 139229 214029
<< labels >>
rlabel metal2 s 938 215988 994 216788 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 57334 215988 57390 216788 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 63038 215988 63094 216788 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 68650 215988 68706 216788 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 74354 215988 74410 216788 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 79966 215988 80022 216788 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 85578 215988 85634 216788 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 91282 215988 91338 216788 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 96894 215988 96950 216788 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 102598 215988 102654 216788 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 108210 215988 108266 216788 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6550 215988 6606 216788 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 113822 215988 113878 216788 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 119526 215988 119582 216788 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 125138 215988 125194 216788 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 130842 215988 130898 216788 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 136454 215988 136510 216788 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 142066 215988 142122 216788 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 147770 215988 147826 216788 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 153382 215988 153438 216788 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 159086 215988 159142 216788 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 164698 215988 164754 216788 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12162 215988 12218 216788 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 170310 215988 170366 216788 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 176014 215988 176070 216788 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 181626 215988 181682 216788 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 187330 215988 187386 216788 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 192942 215988 192998 216788 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 198554 215988 198610 216788 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 204258 215988 204314 216788 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 209870 215988 209926 216788 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 17866 215988 17922 216788 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 23478 215988 23534 216788 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 29090 215988 29146 216788 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 34794 215988 34850 216788 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 40406 215988 40462 216788 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 46110 215988 46166 216788 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 51722 215988 51778 216788 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2778 215988 2834 216788 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 59266 215988 59322 216788 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 64878 215988 64934 216788 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 70582 215988 70638 216788 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 76194 215988 76250 216788 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 81806 215988 81862 216788 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 87510 215988 87566 216788 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 93122 215988 93178 216788 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 98826 215988 98882 216788 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 104438 215988 104494 216788 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 110050 215988 110106 216788 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 8390 215988 8446 216788 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 115754 215988 115810 216788 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 121366 215988 121422 216788 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 127070 215988 127126 216788 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 132682 215988 132738 216788 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 138294 215988 138350 216788 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 143998 215988 144054 216788 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 149610 215988 149666 216788 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 155314 215988 155370 216788 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 160926 215988 160982 216788 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 166538 215988 166594 216788 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 14094 215988 14150 216788 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 172242 215988 172298 216788 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 177854 215988 177910 216788 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 183558 215988 183614 216788 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 189170 215988 189226 216788 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 194782 215988 194838 216788 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 200486 215988 200542 216788 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 206098 215988 206154 216788 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 211802 215988 211858 216788 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 19706 215988 19762 216788 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 25410 215988 25466 216788 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 31022 215988 31078 216788 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 36634 215988 36690 216788 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 42338 215988 42394 216788 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 47950 215988 48006 216788 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 53654 215988 53710 216788 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4618 215988 4674 216788 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 61106 215988 61162 216788 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 66810 215988 66866 216788 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 72422 215988 72478 216788 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 78126 215988 78182 216788 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 83738 215988 83794 216788 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 89350 215988 89406 216788 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 95054 215988 95110 216788 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 100666 215988 100722 216788 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 106370 215988 106426 216788 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 111982 215988 112038 216788 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 10322 215988 10378 216788 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 117594 215988 117650 216788 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 123298 215988 123354 216788 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 128910 215988 128966 216788 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 134614 215988 134670 216788 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 140226 215988 140282 216788 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 145838 215988 145894 216788 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 151542 215988 151598 216788 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 157154 215988 157210 216788 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 162766 215988 162822 216788 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 168470 215988 168526 216788 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 15934 215988 15990 216788 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 174082 215988 174138 216788 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 179786 215988 179842 216788 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 185398 215988 185454 216788 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 191010 215988 191066 216788 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 196714 215988 196770 216788 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 202326 215988 202382 216788 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 208030 215988 208086 216788 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 213642 215988 213698 216788 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 21638 215988 21694 216788 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 27250 215988 27306 216788 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 32862 215988 32918 216788 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 38566 215988 38622 216788 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 44178 215988 44234 216788 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 49882 215988 49938 216788 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 55494 215988 55550 216788 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 213458 0 213514 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 214378 0 214434 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 187330 0 187386 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 212170 0 212226 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 179970 0 180026 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 182546 0 182602 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 185214 0 185270 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 186502 0 186558 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 187790 0 187846 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 193034 0 193090 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 195610 0 195666 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 196898 0 196954 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 198278 0 198334 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 199566 0 199622 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 200854 0 200910 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 203430 0 203486 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 207386 0 207442 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 208674 0 208730 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 209962 0 210018 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 211342 0 211398 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 134246 0 134302 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 172150 0 172206 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 176014 0 176070 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 188250 0 188306 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 201314 0 201370 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 207846 0 207902 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 213090 0 213146 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 214384 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 214384 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 214384 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 214384 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 214384 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 214384 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 214384 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 214384 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 214644 216788
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32980380
string GDS_FILE /Users/somasz/Documents/GitHub/mpw_6c/caravel_design/caravel_bitcoin_asic/openlane/btc_miner_top/runs/btc_miner_top/results/finishing/btc_miner_top.magic.gds
string GDS_START 1142304
<< end >>

