magic
tech sky130B
magscale 1 2
timestamp 1669952481
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 89162 700816 89168 700868
rect 89220 700856 89226 700868
rect 96614 700856 96620 700868
rect 89220 700828 96620 700856
rect 89220 700816 89226 700828
rect 96614 700816 96620 700828
rect 96672 700816 96678 700868
rect 95878 700748 95884 700800
rect 95936 700788 95942 700800
rect 154114 700788 154120 700800
rect 95936 700760 154120 700788
rect 95936 700748 95942 700760
rect 154114 700748 154120 700760
rect 154172 700748 154178 700800
rect 24302 700680 24308 700732
rect 24360 700720 24366 700732
rect 100754 700720 100760 700732
rect 24360 700692 100760 700720
rect 24360 700680 24366 700692
rect 100754 700680 100760 700692
rect 100812 700680 100818 700732
rect 8110 700612 8116 700664
rect 8168 700652 8174 700664
rect 99374 700652 99380 700664
rect 8168 700624 99380 700652
rect 8168 700612 8174 700624
rect 99374 700612 99380 700624
rect 99432 700612 99438 700664
rect 87046 700544 87052 700596
rect 87104 700584 87110 700596
rect 283834 700584 283840 700596
rect 87104 700556 283840 700584
rect 87104 700544 87110 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 84194 700476 84200 700528
rect 84252 700516 84258 700528
rect 348786 700516 348792 700528
rect 84252 700488 348792 700516
rect 84252 700476 84258 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 80054 700408 80060 700460
rect 80112 700448 80118 700460
rect 413646 700448 413652 700460
rect 80112 700420 413652 700448
rect 80112 700408 80118 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 77294 700340 77300 700392
rect 77352 700380 77358 700392
rect 478506 700380 478512 700392
rect 77352 700352 478512 700380
rect 77352 700340 77358 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 74534 700272 74540 700324
rect 74592 700312 74598 700324
rect 543458 700312 543464 700324
rect 74592 700284 543464 700312
rect 74592 700272 74598 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 72970 699660 72976 699712
rect 73028 699700 73034 699712
rect 76558 699700 76564 699712
rect 73028 699672 76564 699700
rect 73028 699660 73034 699672
rect 76558 699660 76564 699672
rect 76616 699660 76622 699712
rect 217318 699660 217324 699712
rect 217376 699700 217382 699712
rect 218974 699700 218980 699712
rect 217376 699672 218980 699700
rect 217376 699660 217382 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 95234 698912 95240 698964
rect 95292 698952 95298 698964
rect 105446 698952 105452 698964
rect 95292 698924 105452 698952
rect 95292 698912 95298 698924
rect 105446 698912 105452 698924
rect 105504 698912 105510 698964
rect 72418 696940 72424 696992
rect 72476 696980 72482 696992
rect 580166 696980 580172 696992
rect 72476 696952 580172 696980
rect 72476 696940 72482 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 92566 696192 92572 696244
rect 92624 696232 92630 696244
rect 137830 696232 137836 696244
rect 92624 696204 137836 696232
rect 92624 696192 92630 696204
rect 137830 696192 137836 696204
rect 137888 696192 137894 696244
rect 85574 693404 85580 693456
rect 85632 693444 85638 693456
rect 267642 693444 267648 693456
rect 85632 693416 267648 693444
rect 85632 693404 85638 693416
rect 267642 693404 267648 693416
rect 267700 693404 267706 693456
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 102134 683244 102140 683256
rect 3476 683216 102140 683244
rect 3476 683204 3482 683216
rect 102134 683204 102140 683216
rect 102192 683204 102198 683256
rect 70486 683136 70492 683188
rect 70544 683176 70550 683188
rect 580166 683176 580172 683188
rect 70544 683148 580172 683176
rect 70544 683136 70550 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 103606 670732 103612 670744
rect 3568 670704 103612 670732
rect 3568 670692 3574 670704
rect 103606 670692 103612 670704
rect 103664 670692 103670 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 102226 656928 102232 656940
rect 3476 656900 102232 656928
rect 3476 656888 3482 656900
rect 102226 656888 102232 656900
rect 102284 656888 102290 656940
rect 66254 643084 66260 643136
rect 66312 643124 66318 643136
rect 580166 643124 580172 643136
rect 66312 643096 580172 643124
rect 66312 643084 66318 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 104894 632108 104900 632120
rect 3476 632080 104900 632108
rect 3476 632068 3482 632080
rect 104894 632068 104900 632080
rect 104952 632068 104958 632120
rect 67634 630640 67640 630692
rect 67692 630680 67698 630692
rect 579982 630680 579988 630692
rect 67692 630652 579988 630680
rect 67692 630640 67698 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 107654 618304 107660 618316
rect 3200 618276 107660 618304
rect 3200 618264 3206 618276
rect 107654 618264 107660 618276
rect 107712 618264 107718 618316
rect 64966 616836 64972 616888
rect 65024 616876 65030 616888
rect 580166 616876 580172 616888
rect 65024 616848 580172 616876
rect 65024 616836 65030 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 106274 605860 106280 605872
rect 3292 605832 106280 605860
rect 3292 605820 3298 605832
rect 106274 605820 106280 605832
rect 106332 605820 106338 605872
rect 63494 590656 63500 590708
rect 63552 590696 63558 590708
rect 580166 590696 580172 590708
rect 63552 590668 580172 590696
rect 63552 590656 63558 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 107746 579680 107752 579692
rect 3384 579652 107752 579680
rect 3384 579640 3390 579652
rect 107746 579640 107752 579652
rect 107804 579640 107810 579692
rect 63586 576852 63592 576904
rect 63644 576892 63650 576904
rect 580166 576892 580172 576904
rect 63644 576864 580172 576892
rect 63644 576852 63650 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 110414 565876 110420 565888
rect 3476 565848 110420 565876
rect 3476 565836 3482 565848
rect 110414 565836 110420 565848
rect 110472 565836 110478 565888
rect 62114 563048 62120 563100
rect 62172 563088 62178 563100
rect 580166 563088 580172 563100
rect 62172 563060 580172 563088
rect 62172 563048 62178 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 109126 553432 109132 553444
rect 3476 553404 109132 553432
rect 3476 553392 3482 553404
rect 109126 553392 109132 553404
rect 109184 553392 109190 553444
rect 59446 536800 59452 536852
rect 59504 536840 59510 536852
rect 579890 536840 579896 536852
rect 59504 536812 579896 536840
rect 59504 536800 59510 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 111794 527184 111800 527196
rect 3476 527156 111800 527184
rect 3476 527144 3482 527156
rect 111794 527144 111800 527156
rect 111852 527144 111858 527196
rect 60734 524424 60740 524476
rect 60792 524464 60798 524476
rect 580166 524464 580172 524476
rect 60792 524436 580172 524464
rect 60792 524424 60798 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 113174 514808 113180 514820
rect 3476 514780 113180 514808
rect 3476 514768 3482 514780
rect 113174 514768 113180 514780
rect 113232 514768 113238 514820
rect 57974 510620 57980 510672
rect 58032 510660 58038 510672
rect 580166 510660 580172 510672
rect 58032 510632 580172 510660
rect 58032 510620 58038 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 113266 501004 113272 501016
rect 3108 500976 113272 501004
rect 3108 500964 3114 500976
rect 113266 500964 113272 500976
rect 113324 500964 113330 501016
rect 40034 496068 40040 496120
rect 40092 496108 40098 496120
rect 98086 496108 98092 496120
rect 40092 496080 98092 496108
rect 40092 496068 40098 496080
rect 98086 496068 98092 496080
rect 98144 496068 98150 496120
rect 88334 494708 88340 494760
rect 88392 494748 88398 494760
rect 234614 494748 234620 494760
rect 88392 494720 234620 494748
rect 88392 494708 88398 494720
rect 234614 494708 234620 494720
rect 234672 494708 234678 494760
rect 56594 484372 56600 484424
rect 56652 484412 56658 484424
rect 580166 484412 580172 484424
rect 56652 484384 580172 484412
rect 56652 484372 56658 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 114646 474756 114652 474768
rect 3476 474728 114652 474756
rect 3476 474716 3482 474728
rect 114646 474716 114652 474728
rect 114704 474716 114710 474768
rect 58066 470568 58072 470620
rect 58124 470608 58130 470620
rect 580166 470608 580172 470620
rect 58124 470580 580172 470608
rect 58124 470568 58130 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 117314 462380 117320 462392
rect 3292 462352 117320 462380
rect 3292 462340 3298 462352
rect 117314 462340 117320 462352
rect 117372 462340 117378 462392
rect 55214 456764 55220 456816
rect 55272 456804 55278 456816
rect 580166 456804 580172 456816
rect 55272 456776 580172 456804
rect 55272 456764 55278 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 115934 448576 115940 448588
rect 3200 448548 115940 448576
rect 3200 448536 3206 448548
rect 115934 448536 115940 448548
rect 115992 448536 115998 448588
rect 52454 430584 52460 430636
rect 52512 430624 52518 430636
rect 579890 430624 579896 430636
rect 52512 430596 579896 430624
rect 52512 430584 52518 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 35158 422328 35164 422340
rect 3476 422300 35164 422328
rect 3476 422288 3482 422300
rect 35158 422288 35164 422300
rect 35216 422288 35222 422340
rect 53926 418140 53932 418192
rect 53984 418180 53990 418192
rect 580166 418180 580172 418192
rect 53984 418152 580172 418180
rect 53984 418140 53990 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 120166 409884 120172 409896
rect 3200 409856 120172 409884
rect 3200 409844 3206 409856
rect 120166 409844 120172 409856
rect 120224 409844 120230 409896
rect 52546 404336 52552 404388
rect 52604 404376 52610 404388
rect 580166 404376 580172 404388
rect 52604 404348 580172 404376
rect 52604 404336 52610 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 94498 397508 94504 397520
rect 3476 397480 94504 397508
rect 3476 397468 3482 397480
rect 94498 397468 94504 397480
rect 94556 397468 94562 397520
rect 49694 378156 49700 378208
rect 49752 378196 49758 378208
rect 580166 378196 580172 378208
rect 49752 378168 580172 378196
rect 49752 378156 49758 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 121454 371260 121460 371272
rect 3476 371232 121460 371260
rect 3476 371220 3482 371232
rect 121454 371220 121460 371232
rect 121512 371220 121518 371272
rect 51074 364352 51080 364404
rect 51132 364392 51138 364404
rect 579614 364392 579620 364404
rect 51132 364364 579620 364392
rect 51132 364352 51138 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 124214 357456 124220 357468
rect 3200 357428 124220 357456
rect 3200 357416 3206 357428
rect 124214 357416 124220 357428
rect 124272 357416 124278 357468
rect 48406 351908 48412 351960
rect 48464 351948 48470 351960
rect 580166 351948 580172 351960
rect 48464 351920 580172 351948
rect 48464 351908 48470 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 122834 345080 122840 345092
rect 3384 345052 122840 345080
rect 3384 345040 3390 345052
rect 122834 345040 122840 345052
rect 122892 345040 122898 345092
rect 46934 324300 46940 324352
rect 46992 324340 46998 324352
rect 580166 324340 580172 324352
rect 46992 324312 580172 324340
rect 46992 324300 46998 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 124306 318832 124312 318844
rect 3476 318804 124312 318832
rect 3476 318792 3482 318804
rect 124306 318792 124312 318804
rect 124364 318792 124370 318844
rect 47026 311856 47032 311908
rect 47084 311896 47090 311908
rect 579982 311896 579988 311908
rect 47084 311868 579988 311896
rect 47084 311856 47090 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 126974 305028 126980 305040
rect 3292 305000 126980 305028
rect 3292 304988 3298 305000
rect 126974 304988 126980 305000
rect 127032 304988 127038 305040
rect 45554 298120 45560 298172
rect 45612 298160 45618 298172
rect 580166 298160 580172 298172
rect 45612 298132 580172 298160
rect 45612 298120 45618 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 125686 292584 125692 292596
rect 3476 292556 125692 292584
rect 3476 292544 3482 292556
rect 125686 292544 125692 292556
rect 125744 292544 125750 292596
rect 42886 271872 42892 271924
rect 42944 271912 42950 271924
rect 580166 271912 580172 271924
rect 42944 271884 580172 271912
rect 42944 271872 42950 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 128354 266404 128360 266416
rect 3108 266376 128360 266404
rect 3108 266364 3114 266376
rect 128354 266364 128360 266376
rect 128412 266364 128418 266416
rect 44174 258068 44180 258120
rect 44232 258108 44238 258120
rect 580166 258108 580172 258120
rect 44232 258080 580172 258108
rect 44232 258068 44238 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 129734 253960 129740 253972
rect 3476 253932 129740 253960
rect 3476 253920 3482 253932
rect 129734 253920 129740 253932
rect 129792 253920 129798 253972
rect 41414 244264 41420 244316
rect 41472 244304 41478 244316
rect 580166 244304 580172 244316
rect 41472 244276 580172 244304
rect 41472 244264 41478 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 3418 240116 3424 240168
rect 3476 240156 3482 240168
rect 129826 240156 129832 240168
rect 3476 240128 129832 240156
rect 3476 240116 3482 240128
rect 129826 240116 129832 240128
rect 129884 240116 129890 240168
rect 40034 231820 40040 231872
rect 40092 231860 40098 231872
rect 579798 231860 579804 231872
rect 40092 231832 579804 231860
rect 40092 231820 40098 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 41506 218016 41512 218068
rect 41564 218056 41570 218068
rect 579890 218056 579896 218068
rect 41564 218028 579896 218056
rect 41564 218016 41570 218028
rect 579890 218016 579896 218028
rect 579948 218016 579954 218068
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 131206 213976 131212 213988
rect 3200 213948 131212 213976
rect 3200 213936 3206 213948
rect 131206 213936 131212 213948
rect 131264 213936 131270 213988
rect 38654 205640 38660 205692
rect 38712 205680 38718 205692
rect 580166 205680 580172 205692
rect 38712 205652 580172 205680
rect 38712 205640 38718 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 3418 201492 3424 201544
rect 3476 201532 3482 201544
rect 133874 201532 133880 201544
rect 3476 201504 133880 201532
rect 3476 201492 3482 201504
rect 133874 201492 133880 201504
rect 133932 201492 133938 201544
rect 35894 191836 35900 191888
rect 35952 191876 35958 191888
rect 580166 191876 580172 191888
rect 35952 191848 580172 191876
rect 35952 191836 35958 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 3418 187688 3424 187740
rect 3476 187728 3482 187740
rect 132494 187728 132500 187740
rect 3476 187700 132500 187728
rect 3476 187688 3482 187700
rect 132494 187688 132500 187700
rect 132552 187688 132558 187740
rect 37366 178032 37372 178084
rect 37424 178072 37430 178084
rect 580166 178072 580172 178084
rect 37424 178044 580172 178072
rect 37424 178032 37430 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 91094 173136 91100 173188
rect 91152 173176 91158 173188
rect 217318 173176 217324 173188
rect 91152 173148 217324 173176
rect 91152 173136 91158 173148
rect 217318 173136 217324 173148
rect 217376 173136 217382 173188
rect 89714 171776 89720 171828
rect 89772 171816 89778 171828
rect 201494 171816 201500 171828
rect 89772 171788 201500 171816
rect 89772 171776 89778 171788
rect 201494 171776 201500 171788
rect 201552 171776 201558 171828
rect 76558 170348 76564 170400
rect 76616 170388 76622 170400
rect 96706 170388 96712 170400
rect 76616 170360 96712 170388
rect 76616 170348 76622 170360
rect 96706 170348 96712 170360
rect 96764 170348 96770 170400
rect 83182 168988 83188 169040
rect 83240 169028 83246 169040
rect 331214 169028 331220 169040
rect 83240 169000 331220 169028
rect 83240 168988 83246 169000
rect 331214 168988 331220 169000
rect 331272 168988 331278 169040
rect 80146 167628 80152 167680
rect 80204 167668 80210 167680
rect 396718 167668 396724 167680
rect 80204 167640 396724 167668
rect 80204 167628 80210 167640
rect 396718 167628 396724 167640
rect 396776 167628 396782 167680
rect 35986 165588 35992 165640
rect 36044 165628 36050 165640
rect 580166 165628 580172 165640
rect 36044 165600 580172 165628
rect 36044 165588 36050 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 76558 164840 76564 164892
rect 76616 164880 76622 164892
rect 462314 164880 462320 164892
rect 76616 164852 462320 164880
rect 76616 164840 76622 164852
rect 462314 164840 462320 164852
rect 462372 164840 462378 164892
rect 3418 162868 3424 162920
rect 3476 162908 3482 162920
rect 135254 162908 135260 162920
rect 3476 162880 135260 162908
rect 3476 162868 3482 162880
rect 135254 162868 135260 162880
rect 135312 162868 135318 162920
rect 33778 162324 33784 162376
rect 33836 162364 33842 162376
rect 119522 162364 119528 162376
rect 33836 162336 119528 162364
rect 33836 162324 33842 162336
rect 119522 162324 119528 162336
rect 119580 162324 119586 162376
rect 20622 162256 20628 162308
rect 20680 162296 20686 162308
rect 151814 162296 151820 162308
rect 20680 162268 151820 162296
rect 20680 162256 20686 162268
rect 151814 162256 151820 162268
rect 151872 162256 151878 162308
rect 2866 162188 2872 162240
rect 2924 162228 2930 162240
rect 153838 162228 153844 162240
rect 2924 162200 153844 162228
rect 2924 162188 2930 162200
rect 153838 162188 153844 162200
rect 153896 162188 153902 162240
rect 1210 162120 1216 162172
rect 1268 162160 1274 162172
rect 188338 162160 188344 162172
rect 1268 162132 188344 162160
rect 1268 162120 1274 162132
rect 188338 162120 188344 162132
rect 188396 162120 188402 162172
rect 3326 162052 3332 162104
rect 3384 162092 3390 162104
rect 196618 162092 196624 162104
rect 3384 162064 196624 162092
rect 3384 162052 3390 162064
rect 196618 162052 196624 162064
rect 196676 162052 196682 162104
rect 17034 161984 17040 162036
rect 17092 162024 17098 162036
rect 220078 162024 220084 162036
rect 17092 161996 220084 162024
rect 17092 161984 17098 161996
rect 220078 161984 220084 161996
rect 220136 161984 220142 162036
rect 12710 161916 12716 161968
rect 12768 161956 12774 161968
rect 233878 161956 233884 161968
rect 12768 161928 233884 161956
rect 12768 161916 12774 161928
rect 233878 161916 233884 161928
rect 233936 161916 233942 161968
rect 4062 161848 4068 161900
rect 4120 161888 4126 161900
rect 285674 161888 285680 161900
rect 4120 161860 285680 161888
rect 4120 161848 4126 161860
rect 285674 161848 285680 161860
rect 285732 161848 285738 161900
rect 8294 161780 8300 161832
rect 8352 161820 8358 161832
rect 302878 161820 302884 161832
rect 8352 161792 302884 161820
rect 8352 161780 8358 161792
rect 302878 161780 302884 161792
rect 302936 161780 302942 161832
rect 8386 161712 8392 161764
rect 8444 161752 8450 161764
rect 305638 161752 305644 161764
rect 8444 161724 305644 161752
rect 8444 161712 8450 161724
rect 305638 161712 305644 161724
rect 305696 161712 305702 161764
rect 2774 161644 2780 161696
rect 2832 161684 2838 161696
rect 309778 161684 309784 161696
rect 2832 161656 309784 161684
rect 2832 161644 2838 161656
rect 309778 161644 309784 161656
rect 309836 161644 309842 161696
rect 15838 161576 15844 161628
rect 15896 161616 15902 161628
rect 422938 161616 422944 161628
rect 15896 161588 422944 161616
rect 15896 161576 15902 161588
rect 422938 161576 422944 161588
rect 422996 161576 423002 161628
rect 7650 161508 7656 161560
rect 7708 161548 7714 161560
rect 449158 161548 449164 161560
rect 7708 161520 449164 161548
rect 7708 161508 7714 161520
rect 449158 161508 449164 161520
rect 449216 161508 449222 161560
rect 69658 161440 69664 161492
rect 69716 161480 69722 161492
rect 557534 161480 557540 161492
rect 69716 161452 557540 161480
rect 69716 161440 69722 161452
rect 557534 161440 557540 161452
rect 557592 161440 557598 161492
rect 69566 160964 69572 161016
rect 69624 161004 69630 161016
rect 201954 161004 201960 161016
rect 69624 160976 201960 161004
rect 69624 160964 69630 160976
rect 201954 160964 201960 160976
rect 202012 160964 202018 161016
rect 12342 160896 12348 160948
rect 12400 160936 12406 160948
rect 150710 160936 150716 160948
rect 12400 160908 150716 160936
rect 12400 160896 12406 160908
rect 150710 160896 150716 160908
rect 150768 160896 150774 160948
rect 12526 160828 12532 160880
rect 12584 160868 12590 160880
rect 152642 160868 152648 160880
rect 12584 160840 152648 160868
rect 12584 160828 12590 160840
rect 152642 160828 152648 160840
rect 152700 160828 152706 160880
rect 2682 160760 2688 160812
rect 2740 160800 2746 160812
rect 174538 160800 174544 160812
rect 2740 160772 174544 160800
rect 2740 160760 2746 160772
rect 174538 160760 174544 160772
rect 174596 160760 174602 160812
rect 35158 160692 35164 160744
rect 35216 160732 35222 160744
rect 118694 160732 118700 160744
rect 35216 160704 118700 160732
rect 35216 160692 35222 160704
rect 118694 160692 118700 160704
rect 118752 160692 118758 160744
rect 119522 160692 119528 160744
rect 119580 160732 119586 160744
rect 295978 160732 295984 160744
rect 119580 160704 295984 160732
rect 119580 160692 119586 160704
rect 295978 160692 295984 160704
rect 296036 160692 296042 160744
rect 3970 160624 3976 160676
rect 4028 160664 4034 160676
rect 215938 160664 215944 160676
rect 4028 160636 215944 160664
rect 4028 160624 4034 160636
rect 215938 160624 215944 160636
rect 215996 160624 216002 160676
rect 3694 160556 3700 160608
rect 3752 160596 3758 160608
rect 246298 160596 246304 160608
rect 3752 160568 246304 160596
rect 3752 160556 3758 160568
rect 246298 160556 246304 160568
rect 246356 160556 246362 160608
rect 73246 160488 73252 160540
rect 73304 160528 73310 160540
rect 353938 160528 353944 160540
rect 73304 160500 353944 160528
rect 73304 160488 73310 160500
rect 353938 160488 353944 160500
rect 353996 160488 354002 160540
rect 2406 160420 2412 160472
rect 2464 160460 2470 160472
rect 283558 160460 283564 160472
rect 2464 160432 283564 160460
rect 2464 160420 2470 160432
rect 283558 160420 283564 160432
rect 283616 160420 283622 160472
rect 20254 160352 20260 160404
rect 20312 160392 20318 160404
rect 335998 160392 336004 160404
rect 20312 160364 336004 160392
rect 20312 160352 20318 160364
rect 335998 160352 336004 160364
rect 336056 160352 336062 160404
rect 13262 160284 13268 160336
rect 13320 160324 13326 160336
rect 381538 160324 381544 160336
rect 13320 160296 381544 160324
rect 13320 160284 13326 160296
rect 381538 160284 381544 160296
rect 381596 160284 381602 160336
rect 3786 160216 3792 160268
rect 3844 160256 3850 160268
rect 400214 160256 400220 160268
rect 3844 160228 400220 160256
rect 3844 160216 3850 160228
rect 400214 160216 400220 160228
rect 400272 160216 400278 160268
rect 3878 160148 3884 160200
rect 3936 160188 3942 160200
rect 445018 160188 445024 160200
rect 3936 160160 445024 160188
rect 3936 160148 3942 160160
rect 445018 160148 445024 160160
rect 445076 160148 445082 160200
rect 2590 160080 2596 160132
rect 2648 160120 2654 160132
rect 463694 160120 463700 160132
rect 2648 160092 463700 160120
rect 2648 160080 2654 160092
rect 463694 160080 463700 160092
rect 463752 160080 463758 160132
rect 5074 159672 5080 159724
rect 5132 159712 5138 159724
rect 20622 159712 20628 159724
rect 5132 159684 20628 159712
rect 5132 159672 5138 159684
rect 20622 159672 20628 159684
rect 20680 159672 20686 159724
rect 18414 159604 18420 159656
rect 18472 159644 18478 159656
rect 33778 159644 33784 159656
rect 18472 159616 33784 159644
rect 18472 159604 18478 159616
rect 33778 159604 33784 159616
rect 33836 159604 33842 159656
rect 73338 159604 73344 159656
rect 73396 159644 73402 159656
rect 156598 159644 156604 159656
rect 73396 159616 156604 159644
rect 73396 159604 73402 159616
rect 156598 159604 156604 159616
rect 156656 159604 156662 159656
rect 6822 159536 6828 159588
rect 6880 159576 6886 159588
rect 12710 159576 12716 159588
rect 6880 159548 12716 159576
rect 6880 159536 6886 159548
rect 12710 159536 12716 159548
rect 12768 159536 12774 159588
rect 16666 159536 16672 159588
rect 16724 159576 16730 159588
rect 150802 159576 150808 159588
rect 16724 159548 150808 159576
rect 16724 159536 16730 159548
rect 150802 159536 150808 159548
rect 150860 159536 150866 159588
rect 9398 159468 9404 159520
rect 9456 159508 9462 159520
rect 152458 159508 152464 159520
rect 9456 159480 152464 159508
rect 9456 159468 9462 159480
rect 152458 159468 152464 159480
rect 152516 159468 152522 159520
rect 11974 159400 11980 159452
rect 12032 159440 12038 159452
rect 161474 159440 161480 159452
rect 12032 159412 161480 159440
rect 12032 159400 12038 159412
rect 161474 159400 161480 159412
rect 161532 159400 161538 159452
rect 6730 159332 6736 159384
rect 6788 159372 6794 159384
rect 180058 159372 180064 159384
rect 6788 159344 180064 159372
rect 6788 159332 6794 159344
rect 180058 159332 180064 159344
rect 180116 159332 180122 159384
rect 6638 159264 6644 159316
rect 6696 159304 6702 159316
rect 251266 159304 251272 159316
rect 6696 159276 251272 159304
rect 6696 159264 6702 159276
rect 251266 159264 251272 159276
rect 251324 159264 251330 159316
rect 6546 159196 6552 159248
rect 6604 159236 6610 159248
rect 267734 159236 267740 159248
rect 6604 159208 267740 159236
rect 6604 159196 6610 159208
rect 267734 159196 267740 159208
rect 267792 159196 267798 159248
rect 934 159128 940 159180
rect 992 159168 998 159180
rect 300118 159168 300124 159180
rect 992 159140 300124 159168
rect 992 159128 998 159140
rect 300118 159128 300124 159140
rect 300176 159128 300182 159180
rect 69658 159060 69664 159112
rect 69716 159100 69722 159112
rect 386414 159100 386420 159112
rect 69716 159072 386420 159100
rect 69716 159060 69722 159072
rect 386414 159060 386420 159072
rect 386472 159060 386478 159112
rect 18782 158992 18788 159044
rect 18840 159032 18846 159044
rect 341518 159032 341524 159044
rect 18840 159004 341524 159032
rect 18840 158992 18846 159004
rect 341518 158992 341524 159004
rect 341576 158992 341582 159044
rect 14274 158924 14280 158976
rect 14332 158964 14338 158976
rect 373994 158964 374000 158976
rect 14332 158936 374000 158964
rect 14332 158924 14338 158936
rect 373994 158924 374000 158936
rect 374052 158924 374058 158976
rect 2314 158856 2320 158908
rect 2372 158896 2378 158908
rect 8294 158896 8300 158908
rect 2372 158868 8300 158896
rect 2372 158856 2378 158868
rect 8294 158856 8300 158868
rect 8352 158856 8358 158908
rect 12618 158856 12624 158908
rect 12676 158896 12682 158908
rect 388438 158896 388444 158908
rect 12676 158868 388444 158896
rect 12676 158856 12682 158868
rect 388438 158856 388444 158868
rect 388496 158856 388502 158908
rect 1026 158788 1032 158840
rect 1084 158828 1090 158840
rect 2866 158828 2872 158840
rect 1084 158800 2872 158828
rect 1084 158788 1090 158800
rect 2866 158788 2872 158800
rect 2924 158788 2930 158840
rect 5442 158788 5448 158840
rect 5500 158828 5506 158840
rect 385678 158828 385684 158840
rect 5500 158800 385684 158828
rect 5500 158788 5506 158800
rect 385678 158788 385684 158800
rect 385736 158788 385742 158840
rect 1302 158720 1308 158772
rect 1360 158760 1366 158772
rect 2774 158760 2780 158772
rect 1360 158732 2780 158760
rect 1360 158720 1366 158732
rect 2774 158720 2780 158732
rect 2832 158720 2838 158772
rect 5350 158720 5356 158772
rect 5408 158760 5414 158772
rect 421558 158760 421564 158772
rect 5408 158732 421564 158760
rect 5408 158720 5414 158732
rect 421558 158720 421564 158732
rect 421616 158720 421622 158772
rect 94498 158244 94504 158296
rect 94556 158284 94562 158296
rect 119706 158284 119712 158296
rect 94556 158256 119712 158284
rect 94556 158244 94562 158256
rect 119706 158244 119712 158256
rect 119764 158244 119770 158296
rect 20346 158176 20352 158228
rect 20404 158216 20410 158228
rect 73246 158216 73252 158228
rect 20404 158188 73252 158216
rect 20404 158176 20410 158188
rect 73246 158176 73252 158188
rect 73304 158176 73310 158228
rect 78582 158176 78588 158228
rect 78640 158216 78646 158228
rect 155862 158216 155868 158228
rect 78640 158188 155868 158216
rect 78640 158176 78646 158188
rect 155862 158176 155868 158188
rect 155920 158176 155926 158228
rect 6178 158108 6184 158160
rect 6236 158148 6242 158160
rect 69566 158148 69572 158160
rect 6236 158120 69572 158148
rect 6236 158108 6242 158120
rect 69566 158108 69572 158120
rect 69624 158108 69630 158160
rect 73154 158108 73160 158160
rect 73212 158148 73218 158160
rect 191098 158148 191104 158160
rect 73212 158120 191104 158148
rect 73212 158108 73218 158120
rect 191098 158108 191104 158120
rect 191156 158108 191162 158160
rect 9674 158040 9680 158092
rect 9732 158080 9738 158092
rect 151906 158080 151912 158092
rect 9732 158052 151912 158080
rect 9732 158040 9738 158052
rect 151906 158040 151912 158052
rect 151964 158040 151970 158092
rect 5166 157972 5172 158024
rect 5224 158012 5230 158024
rect 154022 158012 154028 158024
rect 5224 157984 154028 158012
rect 5224 157972 5230 157984
rect 154022 157972 154028 157984
rect 154080 157972 154086 158024
rect 1118 157904 1124 157956
rect 1176 157944 1182 157956
rect 8386 157944 8392 157956
rect 1176 157916 8392 157944
rect 1176 157904 1182 157916
rect 8386 157904 8392 157916
rect 8444 157904 8450 157956
rect 9306 157904 9312 157956
rect 9364 157944 9370 157956
rect 238018 157944 238024 157956
rect 9364 157916 238024 157944
rect 9364 157904 9370 157916
rect 238018 157904 238024 157916
rect 238076 157904 238082 157956
rect 13722 157836 13728 157888
rect 13780 157876 13786 157888
rect 331214 157876 331220 157888
rect 13780 157848 331220 157876
rect 13780 157836 13786 157848
rect 331214 157836 331220 157848
rect 331272 157836 331278 157888
rect 17402 157768 17408 157820
rect 17460 157808 17466 157820
rect 345658 157808 345664 157820
rect 17460 157780 345664 157808
rect 17460 157768 17466 157780
rect 345658 157768 345664 157780
rect 345716 157768 345722 157820
rect 17862 157700 17868 157752
rect 17920 157740 17926 157752
rect 355318 157740 355324 157752
rect 17920 157712 355324 157740
rect 17920 157700 17926 157712
rect 355318 157700 355324 157712
rect 355376 157700 355382 157752
rect 7834 157632 7840 157684
rect 7892 157672 7898 157684
rect 349154 157672 349160 157684
rect 7892 157644 349160 157672
rect 7892 157632 7898 157644
rect 349154 157632 349160 157644
rect 349212 157632 349218 157684
rect 10042 157564 10048 157616
rect 10100 157604 10106 157616
rect 367738 157604 367744 157616
rect 10100 157576 367744 157604
rect 10100 157564 10106 157576
rect 367738 157564 367744 157576
rect 367796 157564 367802 157616
rect 15010 157496 15016 157548
rect 15068 157536 15074 157548
rect 391198 157536 391204 157548
rect 15068 157508 391204 157536
rect 15068 157496 15074 157508
rect 391198 157496 391204 157508
rect 391256 157496 391262 157548
rect 12986 157428 12992 157480
rect 13044 157468 13050 157480
rect 417418 157468 417424 157480
rect 13044 157440 417424 157468
rect 13044 157428 13050 157440
rect 417418 157428 417424 157440
rect 417476 157428 417482 157480
rect 9490 157360 9496 157412
rect 9548 157400 9554 157412
rect 454678 157400 454684 157412
rect 9548 157372 454684 157400
rect 9548 157360 9554 157372
rect 454678 157360 454684 157372
rect 454736 157360 454742 157412
rect 201954 157292 201960 157344
rect 202012 157332 202018 157344
rect 208486 157332 208492 157344
rect 202012 157304 208492 157332
rect 202012 157292 202018 157304
rect 208486 157292 208492 157304
rect 208544 157292 208550 157344
rect 41414 156884 41420 156936
rect 41472 156924 41478 156936
rect 42426 156924 42432 156936
rect 41472 156896 42432 156924
rect 41472 156884 41478 156896
rect 42426 156884 42432 156896
rect 42484 156884 42490 156936
rect 52454 156884 52460 156936
rect 52512 156924 52518 156936
rect 53466 156924 53472 156936
rect 52512 156896 53472 156924
rect 52512 156884 52518 156896
rect 53466 156884 53472 156896
rect 53524 156884 53530 156936
rect 57974 156884 57980 156936
rect 58032 156924 58038 156936
rect 58986 156924 58992 156936
rect 58032 156896 58992 156924
rect 58032 156884 58038 156896
rect 58986 156884 58992 156896
rect 59044 156884 59050 156936
rect 96614 156884 96620 156936
rect 96672 156924 96678 156936
rect 97626 156924 97632 156936
rect 96672 156896 97632 156924
rect 96672 156884 96678 156896
rect 97626 156884 97632 156896
rect 97684 156884 97690 156936
rect 113174 156884 113180 156936
rect 113232 156924 113238 156936
rect 114186 156924 114192 156936
rect 113232 156896 114192 156924
rect 113232 156884 113238 156896
rect 114186 156884 114192 156896
rect 114244 156884 114250 156936
rect 129734 156884 129740 156936
rect 129792 156924 129798 156936
rect 130746 156924 130752 156936
rect 129792 156896 130752 156924
rect 129792 156884 129798 156896
rect 130746 156884 130752 156896
rect 130804 156884 130810 156936
rect 191098 156884 191104 156936
rect 191156 156924 191162 156936
rect 323578 156924 323584 156936
rect 191156 156896 323584 156924
rect 191156 156884 191162 156896
rect 323578 156884 323584 156896
rect 323636 156884 323642 156936
rect 19242 156816 19248 156868
rect 19300 156856 19306 156868
rect 73154 156856 73160 156868
rect 19300 156828 73160 156856
rect 19300 156816 19306 156828
rect 73154 156816 73160 156828
rect 73212 156816 73218 156868
rect 79502 156816 79508 156868
rect 79560 156856 79566 156868
rect 79560 156828 81388 156856
rect 79560 156816 79566 156828
rect 5258 156748 5264 156800
rect 5316 156788 5322 156800
rect 69658 156788 69664 156800
rect 5316 156760 69664 156788
rect 5316 156748 5322 156760
rect 69658 156748 69664 156760
rect 69716 156748 69722 156800
rect 70302 156748 70308 156800
rect 70360 156788 70366 156800
rect 72418 156788 72424 156800
rect 70360 156760 72424 156788
rect 70360 156748 70366 156760
rect 72418 156748 72424 156760
rect 72476 156748 72482 156800
rect 75822 156748 75828 156800
rect 75880 156788 75886 156800
rect 75880 156760 81296 156788
rect 75880 156748 75886 156760
rect 7926 156680 7932 156732
rect 7984 156720 7990 156732
rect 78582 156720 78588 156732
rect 7984 156692 78588 156720
rect 7984 156680 7990 156692
rect 78582 156680 78588 156692
rect 78640 156680 78646 156732
rect 80054 156680 80060 156732
rect 80112 156720 80118 156732
rect 81066 156720 81072 156732
rect 80112 156692 81072 156720
rect 80112 156680 80118 156692
rect 81066 156680 81072 156692
rect 81124 156680 81130 156732
rect 3602 156612 3608 156664
rect 3660 156652 3666 156664
rect 73338 156652 73344 156664
rect 3660 156624 73344 156652
rect 3660 156612 3666 156624
rect 73338 156612 73344 156624
rect 73396 156612 73402 156664
rect 81268 156652 81296 156760
rect 81360 156720 81388 156828
rect 86126 156816 86132 156868
rect 86184 156856 86190 156868
rect 299474 156856 299480 156868
rect 86184 156828 299480 156856
rect 86184 156816 86190 156828
rect 299474 156816 299480 156828
rect 299532 156816 299538 156868
rect 82722 156748 82728 156800
rect 82780 156788 82786 156800
rect 364334 156788 364340 156800
rect 82780 156760 364340 156788
rect 82780 156748 82786 156760
rect 364334 156748 364340 156760
rect 364392 156748 364398 156800
rect 429194 156720 429200 156732
rect 81360 156692 429200 156720
rect 429194 156680 429200 156692
rect 429252 156680 429258 156732
rect 494054 156652 494060 156664
rect 81268 156624 494060 156652
rect 494054 156612 494060 156624
rect 494112 156612 494118 156664
rect 10962 156544 10968 156596
rect 11020 156584 11026 156596
rect 152734 156584 152740 156596
rect 11020 156556 152740 156584
rect 11020 156544 11026 156556
rect 152734 156544 152740 156556
rect 152792 156544 152798 156596
rect 16482 156476 16488 156528
rect 16540 156516 16546 156528
rect 160094 156516 160100 156528
rect 16540 156488 160100 156516
rect 16540 156476 16546 156488
rect 160094 156476 160100 156488
rect 160152 156476 160158 156528
rect 17770 156408 17776 156460
rect 17828 156448 17834 156460
rect 192478 156448 192484 156460
rect 17828 156420 192484 156448
rect 17828 156408 17834 156420
rect 192478 156408 192484 156420
rect 192536 156408 192542 156460
rect 10778 156340 10784 156392
rect 10836 156380 10842 156392
rect 192570 156380 192576 156392
rect 10836 156352 192576 156380
rect 10836 156340 10842 156352
rect 192570 156340 192576 156352
rect 192628 156340 192634 156392
rect 20162 156272 20168 156324
rect 20220 156312 20226 156324
rect 202138 156312 202144 156324
rect 20220 156284 202144 156312
rect 20220 156272 20226 156284
rect 202138 156272 202144 156284
rect 202196 156272 202202 156324
rect 12894 156204 12900 156256
rect 12952 156244 12958 156256
rect 199378 156244 199384 156256
rect 12952 156216 199384 156244
rect 12952 156204 12958 156216
rect 199378 156204 199384 156216
rect 199436 156204 199442 156256
rect 19058 156136 19064 156188
rect 19116 156176 19122 156188
rect 206370 156176 206376 156188
rect 19116 156148 206376 156176
rect 19116 156136 19122 156148
rect 206370 156136 206376 156148
rect 206428 156136 206434 156188
rect 12434 156068 12440 156120
rect 12492 156108 12498 156120
rect 206278 156108 206284 156120
rect 12492 156080 206284 156108
rect 12492 156068 12498 156080
rect 206278 156068 206284 156080
rect 206336 156068 206342 156120
rect 2498 156000 2504 156052
rect 2556 156040 2562 156052
rect 290550 156040 290556 156052
rect 2556 156012 290556 156040
rect 2556 156000 2562 156012
rect 290550 156000 290556 156012
rect 290608 156000 290614 156052
rect 10226 155932 10232 155984
rect 10284 155972 10290 155984
rect 13262 155972 13268 155984
rect 10284 155944 13268 155972
rect 10284 155932 10290 155944
rect 13262 155932 13268 155944
rect 13320 155932 13326 155984
rect 13354 155932 13360 155984
rect 13412 155972 13418 155984
rect 368474 155972 368480 155984
rect 13412 155944 368480 155972
rect 13412 155932 13418 155944
rect 368474 155932 368480 155944
rect 368532 155932 368538 155984
rect 10318 155864 10324 155916
rect 10376 155904 10382 155916
rect 143994 155904 144000 155916
rect 10376 155876 144000 155904
rect 10376 155864 10382 155876
rect 143994 155864 144000 155876
rect 144052 155864 144058 155916
rect 4798 155796 4804 155848
rect 4856 155836 4862 155848
rect 147306 155836 147312 155848
rect 4856 155808 147312 155836
rect 4856 155796 4862 155808
rect 147306 155796 147312 155808
rect 147364 155796 147370 155848
rect 16390 155728 16396 155780
rect 16448 155768 16454 155780
rect 164234 155768 164240 155780
rect 16448 155740 164240 155768
rect 16448 155728 16454 155740
rect 164234 155728 164240 155740
rect 164292 155728 164298 155780
rect 15930 155660 15936 155712
rect 15988 155700 15994 155712
rect 18782 155700 18788 155712
rect 15988 155672 18788 155700
rect 15988 155660 15994 155672
rect 18782 155660 18788 155672
rect 18840 155660 18846 155712
rect 21358 155660 21364 155712
rect 21416 155700 21422 155712
rect 427078 155700 427084 155712
rect 21416 155672 427084 155700
rect 21416 155660 21422 155672
rect 427078 155660 427084 155672
rect 427136 155660 427142 155712
rect 13262 155592 13268 155644
rect 13320 155632 13326 155644
rect 18046 155632 18052 155644
rect 13320 155604 18052 155632
rect 13320 155592 13326 155604
rect 18046 155592 18052 155604
rect 18104 155592 18110 155644
rect 20898 155592 20904 155644
rect 20956 155632 20962 155644
rect 529934 155632 529940 155644
rect 20956 155604 529940 155632
rect 20956 155592 20962 155604
rect 529934 155592 529940 155604
rect 529992 155592 529998 155644
rect 11882 155524 11888 155576
rect 11940 155564 11946 155576
rect 23474 155564 23480 155576
rect 11940 155536 23480 155564
rect 11940 155524 11946 155536
rect 23474 155524 23480 155536
rect 23532 155524 23538 155576
rect 94958 155524 94964 155576
rect 95016 155564 95022 155576
rect 95878 155564 95884 155576
rect 95016 155536 95884 155564
rect 95016 155524 95022 155536
rect 95878 155524 95884 155536
rect 95936 155524 95942 155576
rect 150434 155524 150440 155576
rect 150492 155564 150498 155576
rect 154114 155564 154120 155576
rect 150492 155536 154120 155564
rect 150492 155524 150498 155536
rect 154114 155524 154120 155536
rect 154172 155524 154178 155576
rect 13446 155456 13452 155508
rect 13504 155496 13510 155508
rect 28810 155496 28816 155508
rect 13504 155468 28816 155496
rect 13504 155456 13510 155468
rect 28810 155456 28816 155468
rect 28868 155456 28874 155508
rect 95602 155456 95608 155508
rect 95660 155496 95666 155508
rect 140774 155496 140780 155508
rect 95660 155468 140780 155496
rect 95660 155456 95666 155468
rect 140774 155456 140780 155468
rect 140832 155456 140838 155508
rect 12250 155388 12256 155440
rect 12308 155428 12314 155440
rect 94314 155428 94320 155440
rect 12308 155400 94320 155428
rect 12308 155388 12314 155400
rect 94314 155388 94320 155400
rect 94372 155388 94378 155440
rect 95694 155388 95700 155440
rect 95752 155428 95758 155440
rect 156506 155428 156512 155440
rect 95752 155400 156512 155428
rect 95752 155388 95758 155400
rect 156506 155388 156512 155400
rect 156564 155388 156570 155440
rect 7742 155320 7748 155372
rect 7800 155360 7806 155372
rect 12618 155360 12624 155372
rect 7800 155332 12624 155360
rect 7800 155320 7806 155332
rect 12618 155320 12624 155332
rect 12676 155320 12682 155372
rect 35250 155320 35256 155372
rect 35308 155360 35314 155372
rect 151170 155360 151176 155372
rect 35308 155332 151176 155360
rect 35308 155320 35314 155332
rect 151170 155320 151176 155332
rect 151228 155320 151234 155372
rect 18322 155252 18328 155304
rect 18380 155292 18386 155304
rect 137370 155292 137376 155304
rect 18380 155264 137376 155292
rect 18380 155252 18386 155264
rect 137370 155252 137376 155264
rect 137428 155252 137434 155304
rect 150526 155252 150532 155304
rect 150584 155292 150590 155304
rect 156690 155292 156696 155304
rect 150584 155264 156696 155292
rect 150584 155252 150590 155264
rect 156690 155252 156696 155264
rect 156748 155252 156754 155304
rect 163498 155252 163504 155304
rect 163556 155292 163562 155304
rect 287698 155292 287704 155304
rect 163556 155264 287704 155292
rect 163556 155252 163562 155264
rect 287698 155252 287704 155264
rect 287756 155252 287762 155304
rect 34146 155184 34152 155236
rect 34204 155224 34210 155236
rect 153102 155224 153108 155236
rect 34204 155196 153108 155224
rect 34204 155184 34210 155196
rect 153102 155184 153108 155196
rect 153160 155184 153166 155236
rect 155862 155184 155868 155236
rect 155920 155224 155926 155236
rect 337378 155224 337384 155236
rect 155920 155196 337384 155224
rect 155920 155184 155926 155196
rect 337378 155184 337384 155196
rect 337436 155184 337442 155236
rect 18506 155116 18512 155168
rect 18564 155156 18570 155168
rect 140958 155156 140964 155168
rect 18564 155128 140964 155156
rect 18564 155116 18570 155128
rect 140958 155116 140964 155128
rect 141016 155116 141022 155168
rect 12066 155048 12072 155100
rect 12124 155088 12130 155100
rect 138014 155088 138020 155100
rect 12124 155060 138020 155088
rect 12124 155048 12130 155060
rect 138014 155048 138020 155060
rect 138072 155048 138078 155100
rect 14366 154980 14372 155032
rect 14424 155020 14430 155032
rect 142890 155020 142896 155032
rect 14424 154992 142896 155020
rect 14424 154980 14430 154992
rect 142890 154980 142896 154992
rect 142948 154980 142954 155032
rect 17218 154912 17224 154964
rect 17276 154952 17282 154964
rect 146294 154952 146300 154964
rect 17276 154924 146300 154952
rect 17276 154912 17282 154924
rect 146294 154912 146300 154924
rect 146352 154912 146358 154964
rect 143350 154844 143356 154896
rect 143408 154884 143414 154896
rect 184934 154884 184940 154896
rect 143408 154856 184940 154884
rect 143408 154844 143414 154856
rect 184934 154844 184940 154856
rect 184992 154844 184998 154896
rect 26234 154776 26240 154828
rect 26292 154816 26298 154828
rect 31018 154816 31024 154828
rect 26292 154788 31024 154816
rect 26292 154776 26298 154788
rect 31018 154776 31024 154788
rect 31076 154776 31082 154828
rect 140866 154776 140872 154828
rect 140924 154816 140930 154828
rect 171134 154816 171140 154828
rect 140924 154788 171140 154816
rect 140924 154776 140930 154788
rect 171134 154776 171140 154788
rect 171192 154776 171198 154828
rect 14642 154708 14648 154760
rect 14700 154748 14706 154760
rect 27522 154748 27528 154760
rect 14700 154720 27528 154748
rect 14700 154708 14706 154720
rect 27522 154708 27528 154720
rect 27580 154708 27586 154760
rect 137186 154708 137192 154760
rect 137244 154748 137250 154760
rect 152918 154748 152924 154760
rect 137244 154720 152924 154748
rect 137244 154708 137250 154720
rect 152918 154708 152924 154720
rect 152976 154708 152982 154760
rect 9582 154640 9588 154692
rect 9640 154680 9646 154692
rect 12986 154680 12992 154692
rect 9640 154652 12992 154680
rect 9640 154640 9646 154652
rect 12986 154640 12992 154652
rect 13044 154640 13050 154692
rect 16298 154640 16304 154692
rect 16356 154680 16362 154692
rect 22186 154680 22192 154692
rect 16356 154652 22192 154680
rect 16356 154640 16362 154652
rect 22186 154640 22192 154652
rect 22244 154640 22250 154692
rect 30190 154640 30196 154692
rect 30248 154680 30254 154692
rect 96522 154680 96528 154692
rect 30248 154652 96528 154680
rect 30248 154640 30254 154652
rect 96522 154640 96528 154652
rect 96580 154640 96586 154692
rect 146754 154640 146760 154692
rect 146812 154680 146818 154692
rect 151446 154680 151452 154692
rect 146812 154652 151452 154680
rect 146812 154640 146818 154652
rect 151446 154640 151452 154652
rect 151504 154640 151510 154692
rect 152826 154680 152832 154692
rect 151786 154652 152832 154680
rect 8110 154572 8116 154624
rect 8168 154612 8174 154624
rect 9674 154612 9680 154624
rect 8168 154584 9680 154612
rect 8168 154572 8174 154584
rect 9674 154572 9680 154584
rect 9732 154572 9738 154624
rect 10870 154572 10876 154624
rect 10928 154612 10934 154624
rect 26234 154612 26240 154624
rect 10928 154584 26240 154612
rect 10928 154572 10934 154584
rect 26234 154572 26240 154584
rect 26292 154572 26298 154624
rect 28902 154612 28908 154624
rect 26436 154584 28908 154612
rect 8294 154504 8300 154556
rect 8352 154544 8358 154556
rect 12342 154544 12348 154556
rect 8352 154516 12348 154544
rect 8352 154504 8358 154516
rect 12342 154504 12348 154516
rect 12400 154504 12406 154556
rect 19610 154504 19616 154556
rect 19668 154544 19674 154556
rect 26436 154544 26464 154584
rect 28902 154572 28908 154584
rect 28960 154572 28966 154624
rect 35894 154572 35900 154624
rect 35952 154612 35958 154624
rect 36906 154612 36912 154624
rect 35952 154584 36912 154612
rect 35952 154572 35958 154584
rect 36906 154572 36912 154584
rect 36964 154572 36970 154624
rect 140774 154572 140780 154624
rect 140832 154612 140838 154624
rect 151786 154612 151814 154652
rect 152826 154640 152832 154652
rect 152884 154640 152890 154692
rect 140832 154584 142154 154612
rect 140832 154572 140838 154584
rect 19668 154516 26464 154544
rect 142126 154544 142154 154584
rect 143552 154584 151814 154612
rect 143552 154544 143580 154584
rect 142126 154516 143580 154544
rect 19668 154504 19674 154516
rect 8938 154232 8944 154284
rect 8996 154272 9002 154284
rect 145098 154272 145104 154284
rect 8996 154244 145104 154272
rect 8996 154232 9002 154244
rect 145098 154232 145104 154244
rect 145156 154232 145162 154284
rect 10410 154164 10416 154216
rect 10468 154204 10474 154216
rect 35710 154204 35716 154216
rect 10468 154176 35716 154204
rect 10468 154164 10474 154176
rect 35710 154164 35716 154176
rect 35768 154164 35774 154216
rect 94314 154164 94320 154216
rect 94372 154204 94378 154216
rect 150526 154204 150532 154216
rect 94372 154176 150532 154204
rect 94372 154164 94378 154176
rect 150526 154164 150532 154176
rect 150584 154164 150590 154216
rect 9214 154096 9220 154148
rect 9272 154136 9278 154148
rect 10042 154136 10048 154148
rect 9272 154108 10048 154136
rect 9272 154096 9278 154108
rect 10042 154096 10048 154108
rect 10100 154096 10106 154148
rect 12158 154096 12164 154148
rect 12216 154136 12222 154148
rect 30282 154136 30288 154148
rect 12216 154108 30288 154136
rect 12216 154096 12222 154108
rect 30282 154096 30288 154108
rect 30340 154096 30346 154148
rect 34422 154096 34428 154148
rect 34480 154136 34486 154148
rect 95694 154136 95700 154148
rect 34480 154108 95700 154136
rect 34480 154096 34486 154108
rect 95694 154096 95700 154108
rect 95752 154096 95758 154148
rect 153102 154096 153108 154148
rect 153160 154136 153166 154148
rect 164786 154136 164792 154148
rect 153160 154108 164792 154136
rect 153160 154096 153166 154108
rect 164786 154096 164792 154108
rect 164844 154096 164850 154148
rect 30926 154028 30932 154080
rect 30984 154068 30990 154080
rect 95142 154068 95148 154080
rect 30984 154040 95148 154068
rect 30984 154028 30990 154040
rect 95142 154028 95148 154040
rect 95200 154028 95206 154080
rect 96522 154028 96528 154080
rect 96580 154068 96586 154080
rect 143442 154068 143448 154080
rect 96580 154040 143448 154068
rect 96580 154028 96586 154040
rect 143442 154028 143448 154040
rect 143500 154028 143506 154080
rect 160094 154028 160100 154080
rect 160152 154068 160158 154080
rect 195606 154068 195612 154080
rect 160152 154040 195612 154068
rect 160152 154028 160158 154040
rect 195606 154028 195612 154040
rect 195664 154028 195670 154080
rect 290550 154028 290556 154080
rect 290608 154068 290614 154080
rect 317414 154068 317420 154080
rect 290608 154040 317420 154068
rect 290608 154028 290614 154040
rect 317414 154028 317420 154040
rect 317472 154028 317478 154080
rect 35802 153960 35808 154012
rect 35860 154000 35866 154012
rect 137278 154000 137284 154012
rect 35860 153972 137284 154000
rect 35860 153960 35866 153972
rect 137278 153960 137284 153972
rect 137336 153960 137342 154012
rect 138014 153960 138020 154012
rect 138072 154000 138078 154012
rect 151354 154000 151360 154012
rect 138072 153972 151360 154000
rect 138072 153960 138078 153972
rect 151354 153960 151360 153972
rect 151412 153960 151418 154012
rect 156598 153960 156604 154012
rect 156656 154000 156662 154012
rect 208394 154000 208400 154012
rect 156656 153972 208400 154000
rect 156656 153960 156662 153972
rect 208394 153960 208400 153972
rect 208452 153960 208458 154012
rect 208486 153960 208492 154012
rect 208544 154000 208550 154012
rect 292482 154000 292488 154012
rect 208544 153972 292488 154000
rect 208544 153960 208550 153972
rect 292482 153960 292488 153972
rect 292540 153960 292546 154012
rect 23474 153892 23480 153944
rect 23532 153932 23538 153944
rect 32950 153932 32956 153944
rect 23532 153904 32956 153932
rect 23532 153892 23538 153904
rect 32950 153892 32956 153904
rect 33008 153892 33014 153944
rect 33042 153892 33048 153944
rect 33100 153932 33106 153944
rect 150434 153932 150440 153944
rect 33100 153904 150440 153932
rect 33100 153892 33106 153904
rect 150434 153892 150440 153904
rect 150492 153892 150498 153944
rect 156506 153892 156512 153944
rect 156564 153932 156570 153944
rect 359458 153932 359464 153944
rect 156564 153904 359464 153932
rect 156564 153892 156570 153904
rect 359458 153892 359464 153904
rect 359516 153892 359522 153944
rect 8202 153824 8208 153876
rect 8260 153864 8266 153876
rect 17862 153864 17868 153876
rect 8260 153836 17868 153864
rect 8260 153824 8266 153836
rect 17862 153824 17868 153836
rect 17920 153824 17926 153876
rect 18138 153824 18144 153876
rect 18196 153864 18202 153876
rect 34146 153864 34152 153876
rect 18196 153836 34152 153864
rect 18196 153824 18202 153836
rect 34146 153824 34152 153836
rect 34204 153824 34210 153876
rect 35618 153824 35624 153876
rect 35676 153864 35682 153876
rect 409138 153864 409144 153876
rect 35676 153836 409144 153864
rect 35676 153824 35682 153836
rect 409138 153824 409144 153836
rect 409196 153824 409202 153876
rect 427078 153824 427084 153876
rect 427136 153864 427142 153876
rect 485038 153864 485044 153876
rect 427136 153836 485044 153864
rect 427136 153824 427142 153836
rect 485038 153824 485044 153836
rect 485096 153824 485102 153876
rect 7558 153756 7564 153808
rect 7616 153796 7622 153808
rect 141786 153796 141792 153808
rect 7616 153768 141792 153796
rect 7616 153756 7622 153768
rect 141786 153756 141792 153768
rect 141844 153756 141850 153808
rect 3234 153688 3240 153740
rect 3292 153728 3298 153740
rect 138474 153728 138480 153740
rect 3292 153700 138480 153728
rect 3292 153688 3298 153700
rect 138474 153688 138480 153700
rect 138532 153688 138538 153740
rect 17678 153620 17684 153672
rect 17736 153660 17742 153672
rect 156598 153660 156604 153672
rect 17736 153632 156604 153660
rect 17736 153620 17742 153632
rect 156598 153620 156604 153632
rect 156656 153620 156662 153672
rect 17494 153552 17500 153604
rect 17552 153592 17558 153604
rect 427078 153592 427084 153604
rect 17552 153564 427084 153592
rect 17552 153552 17558 153564
rect 427078 153552 427084 153564
rect 427136 153552 427142 153604
rect 17586 153484 17592 153536
rect 17644 153524 17650 153536
rect 431218 153524 431224 153536
rect 17644 153496 431224 153524
rect 17644 153484 17650 153496
rect 431218 153484 431224 153496
rect 431276 153484 431282 153536
rect 23198 153416 23204 153468
rect 23256 153456 23262 153468
rect 34974 153456 34980 153468
rect 23256 153428 34980 153456
rect 23256 153416 23262 153428
rect 34974 153416 34980 153428
rect 35032 153416 35038 153468
rect 137094 153416 137100 153468
rect 137152 153456 137158 153468
rect 578878 153456 578884 153468
rect 137152 153428 578884 153456
rect 137152 153416 137158 153428
rect 578878 153416 578884 153428
rect 578936 153416 578942 153468
rect 18782 153348 18788 153400
rect 18840 153388 18846 153400
rect 462958 153388 462964 153400
rect 18840 153360 462964 153388
rect 18840 153348 18846 153360
rect 462958 153348 462964 153360
rect 463016 153348 463022 153400
rect 2222 153280 2228 153332
rect 2280 153320 2286 153332
rect 7650 153320 7656 153332
rect 2280 153292 7656 153320
rect 2280 153280 2286 153292
rect 7650 153280 7656 153292
rect 7708 153280 7714 153332
rect 18690 153280 18696 153332
rect 18748 153320 18754 153332
rect 489914 153320 489920 153332
rect 18748 153292 489920 153320
rect 18748 153280 18754 153292
rect 489914 153280 489920 153292
rect 489972 153280 489978 153332
rect 6454 153212 6460 153264
rect 6512 153252 6518 153264
rect 9398 153252 9404 153264
rect 6512 153224 9404 153252
rect 6512 153212 6518 153224
rect 9398 153212 9404 153224
rect 9456 153212 9462 153264
rect 17862 153212 17868 153264
rect 17920 153252 17926 153264
rect 525794 153252 525800 153264
rect 17920 153224 525800 153252
rect 17920 153212 17926 153224
rect 525794 153212 525800 153224
rect 525852 153212 525858 153264
rect 842 153144 848 153196
rect 900 153184 906 153196
rect 3326 153184 3332 153196
rect 900 153156 3332 153184
rect 900 153144 906 153156
rect 3326 153144 3332 153156
rect 3384 153144 3390 153196
rect 15102 153144 15108 153196
rect 15160 153184 15166 153196
rect 15838 153184 15844 153196
rect 15160 153156 15844 153184
rect 15160 153144 15166 153156
rect 15838 153144 15844 153156
rect 15896 153144 15902 153196
rect 17126 153144 17132 153196
rect 17184 153184 17190 153196
rect 20346 153184 20352 153196
rect 17184 153156 20352 153184
rect 17184 153144 17190 153156
rect 20346 153144 20352 153156
rect 20404 153144 20410 153196
rect 27522 153144 27528 153196
rect 27580 153184 27586 153196
rect 30926 153184 30932 153196
rect 27580 153156 30932 153184
rect 27580 153144 27586 153156
rect 30926 153144 30932 153156
rect 30984 153144 30990 153196
rect 31018 153144 31024 153196
rect 31076 153184 31082 153196
rect 35802 153184 35808 153196
rect 31076 153156 35808 153184
rect 31076 153144 31082 153156
rect 35802 153144 35808 153156
rect 35860 153144 35866 153196
rect 140866 153184 140872 153196
rect 35912 153156 140872 153184
rect 19886 153076 19892 153128
rect 19944 153116 19950 153128
rect 19944 153088 26234 153116
rect 19944 153076 19950 153088
rect 26206 153048 26234 153088
rect 28810 153076 28816 153128
rect 28868 153116 28874 153128
rect 33042 153116 33048 153128
rect 28868 153088 33048 153116
rect 28868 153076 28874 153088
rect 33042 153076 33048 153088
rect 33100 153076 33106 153128
rect 35912 153116 35940 153156
rect 140866 153144 140872 153156
rect 140924 153144 140930 153196
rect 137186 153116 137192 153128
rect 35636 153088 35940 153116
rect 41386 153088 137192 153116
rect 30190 153048 30196 153060
rect 26206 153020 30196 153048
rect 30190 153008 30196 153020
rect 30248 153008 30254 153060
rect 16022 152940 16028 152992
rect 16080 152980 16086 152992
rect 20622 152980 20628 152992
rect 16080 152952 20628 152980
rect 16080 152940 16086 152952
rect 20622 152940 20628 152952
rect 20680 152940 20686 152992
rect 30282 152940 30288 152992
rect 30340 152980 30346 152992
rect 35636 152980 35664 153088
rect 35710 153008 35716 153060
rect 35768 153048 35774 153060
rect 41386 153048 41414 153088
rect 137186 153076 137192 153088
rect 137244 153076 137250 153128
rect 137278 153076 137284 153128
rect 137336 153116 137342 153128
rect 146754 153116 146760 153128
rect 137336 153088 146760 153116
rect 137336 153076 137342 153088
rect 146754 153076 146760 153088
rect 146812 153076 146818 153128
rect 95602 153048 95608 153060
rect 35768 153020 41414 153048
rect 45526 153020 95608 153048
rect 35768 153008 35774 153020
rect 30340 152952 35664 152980
rect 30340 152940 30346 152952
rect 16206 152872 16212 152924
rect 16264 152912 16270 152924
rect 21358 152912 21364 152924
rect 16264 152884 21364 152912
rect 16264 152872 16270 152884
rect 21358 152872 21364 152884
rect 21416 152872 21422 152924
rect 32950 152872 32956 152924
rect 33008 152912 33014 152924
rect 45526 152912 45554 153020
rect 95602 153008 95608 153020
rect 95660 153008 95666 153060
rect 33008 152884 45554 152912
rect 33008 152872 33014 152884
rect 14918 152736 14924 152788
rect 14976 152776 14982 152788
rect 20898 152776 20904 152788
rect 14976 152748 20904 152776
rect 14976 152736 14982 152748
rect 20898 152736 20904 152748
rect 20956 152736 20962 152788
rect 143442 152668 143448 152720
rect 143500 152708 143506 152720
rect 151998 152708 152004 152720
rect 143500 152680 152004 152708
rect 143500 152668 143506 152680
rect 151998 152668 152004 152680
rect 152056 152668 152062 152720
rect 164786 152668 164792 152720
rect 164844 152708 164850 152720
rect 175274 152708 175280 152720
rect 164844 152680 175280 152708
rect 164844 152668 164850 152680
rect 175274 152668 175280 152680
rect 175332 152668 175338 152720
rect 8018 152600 8024 152652
rect 8076 152640 8082 152652
rect 17402 152640 17408 152652
rect 8076 152612 17408 152640
rect 8076 152600 8082 152612
rect 17402 152600 17408 152612
rect 17460 152600 17466 152652
rect 150526 152600 150532 152652
rect 150584 152640 150590 152652
rect 166258 152640 166264 152652
rect 150584 152612 166264 152640
rect 150584 152600 150590 152612
rect 166258 152600 166264 152612
rect 166316 152600 166322 152652
rect 4982 152532 4988 152584
rect 5040 152572 5046 152584
rect 16666 152572 16672 152584
rect 5040 152544 16672 152572
rect 5040 152532 5046 152544
rect 16666 152532 16672 152544
rect 16724 152532 16730 152584
rect 150434 152532 150440 152584
rect 150492 152572 150498 152584
rect 178034 152572 178040 152584
rect 150492 152544 178040 152572
rect 150492 152532 150498 152544
rect 178034 152532 178040 152544
rect 178092 152532 178098 152584
rect 4890 152464 4896 152516
rect 4948 152504 4954 152516
rect 12526 152504 12532 152516
rect 4948 152476 12532 152504
rect 4948 152464 4954 152476
rect 12526 152464 12532 152476
rect 12584 152464 12590 152516
rect 15746 152464 15752 152516
rect 15804 152504 15810 152516
rect 34422 152504 34428 152516
rect 15804 152476 34428 152504
rect 15804 152464 15810 152476
rect 34422 152464 34428 152476
rect 34480 152464 34486 152516
rect 35342 152464 35348 152516
rect 35400 152504 35406 152516
rect 150986 152504 150992 152516
rect 35400 152476 150992 152504
rect 35400 152464 35406 152476
rect 150986 152464 150992 152476
rect 151044 152464 151050 152516
rect 156690 152464 156696 152516
rect 156748 152504 156754 152516
rect 323026 152504 323032 152516
rect 156748 152476 323032 152504
rect 156748 152464 156754 152476
rect 323026 152464 323032 152476
rect 323084 152464 323090 152516
rect 359458 152464 359464 152516
rect 359516 152504 359522 152516
rect 406378 152504 406384 152516
rect 359516 152476 406384 152504
rect 359516 152464 359522 152476
rect 406378 152464 406384 152476
rect 406436 152464 406442 152516
rect 485038 152464 485044 152516
rect 485096 152504 485102 152516
rect 516778 152504 516784 152516
rect 485096 152476 516784 152504
rect 485096 152464 485102 152476
rect 516778 152464 516784 152476
rect 516836 152464 516842 152516
rect 18874 152260 18880 152312
rect 18932 152300 18938 152312
rect 467098 152300 467104 152312
rect 18932 152272 467104 152300
rect 18932 152260 18938 152272
rect 467098 152260 467104 152272
rect 467156 152260 467162 152312
rect 12986 152192 12992 152244
rect 13044 152232 13050 152244
rect 139578 152232 139584 152244
rect 13044 152204 139584 152232
rect 13044 152192 13050 152204
rect 139578 152192 139584 152204
rect 139636 152192 139642 152244
rect 3418 152124 3424 152176
rect 3476 152164 3482 152176
rect 136266 152164 136272 152176
rect 3476 152136 136272 152164
rect 3476 152124 3482 152136
rect 136266 152124 136272 152136
rect 136324 152124 136330 152176
rect 18598 152056 18604 152108
rect 18656 152096 18662 152108
rect 363598 152096 363604 152108
rect 18656 152068 363604 152096
rect 18656 152056 18662 152068
rect 363598 152056 363604 152068
rect 363656 152056 363662 152108
rect 11790 151988 11796 152040
rect 11848 152028 11854 152040
rect 18138 152028 18144 152040
rect 11848 152000 18144 152028
rect 11848 151988 11854 152000
rect 18138 151988 18144 152000
rect 18196 151988 18202 152040
rect 18966 151988 18972 152040
rect 19024 152028 19030 152040
rect 453298 152028 453304 152040
rect 19024 152000 453304 152028
rect 19024 151988 19030 152000
rect 453298 151988 453304 152000
rect 453356 151988 453362 152040
rect 11698 151920 11704 151972
rect 11756 151960 11762 151972
rect 18414 151960 18420 151972
rect 11756 151932 18420 151960
rect 11756 151920 11762 151932
rect 18414 151920 18420 151932
rect 18472 151920 18478 151972
rect 19978 151920 19984 151972
rect 20036 151960 20042 151972
rect 458818 151960 458824 151972
rect 20036 151932 458824 151960
rect 20036 151920 20042 151932
rect 458818 151920 458824 151932
rect 458876 151920 458882 151972
rect 10686 151852 10692 151904
rect 10744 151892 10750 151904
rect 19886 151892 19892 151904
rect 10744 151864 19892 151892
rect 10744 151852 10750 151864
rect 19886 151852 19892 151864
rect 19944 151852 19950 151904
rect 20070 151852 20076 151904
rect 20128 151892 20134 151904
rect 460198 151892 460204 151904
rect 20128 151864 460204 151892
rect 20128 151852 20134 151864
rect 460198 151852 460204 151864
rect 460256 151852 460262 151904
rect 18230 151824 18236 151836
rect 16592 151796 18236 151824
rect 13170 151716 13176 151768
rect 13228 151756 13234 151768
rect 16592 151756 16620 151796
rect 18230 151784 18236 151796
rect 18288 151784 18294 151836
rect 13228 151728 16620 151756
rect 13228 151716 13234 151728
rect 317414 151716 317420 151768
rect 317472 151756 317478 151768
rect 327718 151756 327724 151768
rect 317472 151728 327724 151756
rect 317472 151716 317478 151728
rect 327718 151716 327724 151728
rect 327776 151716 327782 151768
rect 292482 151648 292488 151700
rect 292540 151688 292546 151700
rect 319438 151688 319444 151700
rect 292540 151660 319444 151688
rect 292540 151648 292546 151660
rect 319438 151648 319444 151660
rect 319496 151648 319502 151700
rect 323578 151648 323584 151700
rect 323636 151688 323642 151700
rect 377398 151688 377404 151700
rect 323636 151660 377404 151688
rect 323636 151648 323642 151660
rect 377398 151648 377404 151660
rect 377456 151648 377462 151700
rect 150894 151580 150900 151632
rect 150952 151620 150958 151632
rect 182174 151620 182180 151632
rect 150952 151592 182180 151620
rect 150952 151580 150958 151592
rect 182174 151580 182180 151592
rect 182232 151580 182238 151632
rect 206370 151580 206376 151632
rect 206428 151620 206434 151632
rect 324406 151620 324412 151632
rect 206428 151592 324412 151620
rect 206428 151580 206434 151592
rect 324406 151580 324412 151592
rect 324464 151580 324470 151632
rect 337378 151580 337384 151632
rect 337436 151620 337442 151632
rect 403618 151620 403624 151632
rect 337436 151592 403624 151620
rect 337436 151580 337442 151592
rect 403618 151580 403624 151592
rect 403676 151580 403682 151632
rect 152918 151512 152924 151564
rect 152976 151552 152982 151564
rect 193214 151552 193220 151564
rect 152976 151524 193220 151552
rect 152976 151512 152982 151524
rect 193214 151512 193220 151524
rect 193272 151512 193278 151564
rect 195606 151512 195612 151564
rect 195664 151552 195670 151564
rect 338114 151552 338120 151564
rect 195664 151524 338120 151552
rect 195664 151512 195670 151524
rect 338114 151512 338120 151524
rect 338172 151512 338178 151564
rect 152826 151444 152832 151496
rect 152884 151484 152890 151496
rect 207014 151484 207020 151496
rect 152884 151456 207020 151484
rect 152884 151444 152890 151456
rect 207014 151444 207020 151456
rect 207072 151444 207078 151496
rect 208394 151444 208400 151496
rect 208452 151484 208458 151496
rect 292666 151484 292672 151496
rect 208452 151456 292672 151484
rect 208452 151444 208458 151456
rect 292666 151444 292672 151456
rect 292724 151444 292730 151496
rect 323026 151444 323032 151496
rect 323084 151484 323090 151496
rect 476758 151484 476764 151496
rect 323084 151456 476764 151484
rect 323084 151444 323090 151456
rect 476758 151444 476764 151456
rect 476816 151444 476822 151496
rect 151354 151376 151360 151428
rect 151412 151416 151418 151428
rect 189074 151416 189080 151428
rect 151412 151388 189080 151416
rect 151412 151376 151418 151388
rect 189074 151376 189080 151388
rect 189132 151376 189138 151428
rect 192570 151376 192576 151428
rect 192628 151416 192634 151428
rect 356698 151416 356704 151428
rect 192628 151388 356704 151416
rect 192628 151376 192634 151388
rect 356698 151376 356704 151388
rect 356756 151376 356762 151428
rect 151998 151308 152004 151360
rect 152056 151348 152062 151360
rect 202874 151348 202880 151360
rect 152056 151320 202880 151348
rect 152056 151308 152062 151320
rect 202874 151308 202880 151320
rect 202932 151308 202938 151360
rect 206278 151308 206284 151360
rect 206336 151348 206342 151360
rect 394694 151348 394700 151360
rect 206336 151320 394700 151348
rect 206336 151308 206342 151320
rect 394694 151308 394700 151320
rect 394752 151308 394758 151360
rect 152090 151240 152096 151292
rect 152148 151280 152154 151292
rect 200114 151280 200120 151292
rect 152148 151252 200120 151280
rect 152148 151240 152154 151252
rect 200114 151240 200120 151252
rect 200172 151240 200178 151292
rect 202138 151240 202144 151292
rect 202196 151280 202202 151292
rect 399478 151280 399484 151292
rect 202196 151252 399484 151280
rect 202196 151240 202202 151252
rect 399478 151240 399484 151252
rect 399536 151240 399542 151292
rect 422938 151240 422944 151292
rect 422996 151280 423002 151292
rect 435358 151280 435364 151292
rect 422996 151252 435364 151280
rect 422996 151240 423002 151252
rect 435358 151240 435364 151252
rect 435416 151240 435422 151292
rect 151446 151172 151452 151224
rect 151504 151212 151510 151224
rect 195974 151212 195980 151224
rect 151504 151184 195980 151212
rect 151504 151172 151510 151184
rect 195974 151172 195980 151184
rect 196032 151172 196038 151224
rect 199378 151172 199384 151224
rect 199436 151212 199442 151224
rect 503714 151212 503720 151224
rect 199436 151184 503720 151212
rect 199436 151172 199442 151184
rect 503714 151172 503720 151184
rect 503772 151172 503778 151224
rect 151262 151104 151268 151156
rect 151320 151144 151326 151156
rect 491938 151144 491944 151156
rect 151320 151116 491944 151144
rect 151320 151104 151326 151116
rect 491938 151104 491944 151116
rect 491996 151104 492002 151156
rect 16114 151036 16120 151088
rect 16172 151076 16178 151088
rect 19794 151076 19800 151088
rect 16172 151048 19800 151076
rect 16172 151036 16178 151048
rect 19794 151036 19800 151048
rect 19852 151036 19858 151088
rect 150986 151036 150992 151088
rect 151044 151076 151050 151088
rect 561674 151076 561680 151088
rect 151044 151048 561680 151076
rect 151044 151036 151050 151048
rect 561674 151036 561680 151048
rect 561732 151036 561738 151088
rect 10594 150560 10600 150612
rect 10652 150600 10658 150612
rect 15930 150600 15936 150612
rect 10652 150572 15936 150600
rect 10652 150560 10658 150572
rect 15930 150560 15936 150572
rect 15988 150560 15994 150612
rect 9030 150492 9036 150544
rect 9088 150532 9094 150544
rect 11974 150532 11980 150544
rect 9088 150504 11980 150532
rect 9088 150492 9094 150504
rect 11974 150492 11980 150504
rect 12032 150492 12038 150544
rect 17310 150492 17316 150544
rect 17368 150532 17374 150544
rect 19610 150532 19616 150544
rect 17368 150504 19616 150532
rect 17368 150492 17374 150504
rect 19610 150492 19616 150504
rect 19668 150492 19674 150544
rect 192478 150492 192484 150544
rect 192536 150532 192542 150544
rect 197354 150532 197360 150544
rect 192536 150504 197360 150532
rect 192536 150492 192542 150504
rect 197354 150492 197360 150504
rect 197412 150492 197418 150544
rect 7650 150424 7656 150476
rect 7708 150464 7714 150476
rect 9122 150464 9128 150476
rect 7708 150436 9128 150464
rect 7708 150424 7714 150436
rect 9122 150424 9128 150436
rect 9180 150424 9186 150476
rect 9306 150424 9312 150476
rect 9364 150464 9370 150476
rect 12894 150464 12900 150476
rect 9364 150436 12900 150464
rect 9364 150424 9370 150436
rect 12894 150424 12900 150436
rect 12952 150424 12958 150476
rect 13078 150424 13084 150476
rect 13136 150464 13142 150476
rect 14458 150464 14464 150476
rect 13136 150436 14464 150464
rect 13136 150424 13142 150436
rect 14458 150424 14464 150436
rect 14516 150424 14522 150476
rect 17402 150424 17408 150476
rect 17460 150464 17466 150476
rect 19702 150464 19708 150476
rect 17460 150436 19708 150464
rect 17460 150424 17466 150436
rect 19702 150424 19708 150436
rect 19760 150424 19766 150476
rect 196618 150424 196624 150476
rect 196676 150464 196682 150476
rect 201494 150464 201500 150476
rect 196676 150436 201500 150464
rect 196676 150424 196682 150436
rect 201494 150424 201500 150436
rect 201552 150424 201558 150476
rect 355318 150424 355324 150476
rect 355376 150464 355382 150476
rect 359458 150464 359464 150476
rect 355376 150436 359464 150464
rect 355376 150424 355382 150436
rect 359458 150424 359464 150436
rect 359516 150424 359522 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 18322 150396 18328 150408
rect 3476 150368 18328 150396
rect 3476 150356 3482 150368
rect 18322 150356 18328 150368
rect 18380 150356 18386 150408
rect 154114 149812 154120 149864
rect 154172 149852 154178 149864
rect 278038 149852 278044 149864
rect 154172 149824 278044 149852
rect 154172 149812 154178 149824
rect 278038 149812 278044 149824
rect 278096 149812 278102 149864
rect 154022 149744 154028 149796
rect 154080 149784 154086 149796
rect 313918 149784 313924 149796
rect 154080 149756 313924 149784
rect 154080 149744 154086 149756
rect 313918 149744 313924 149756
rect 313976 149744 313982 149796
rect 15930 149676 15936 149728
rect 15988 149716 15994 149728
rect 17034 149716 17040 149728
rect 15988 149688 17040 149716
rect 15988 149676 15994 149688
rect 17034 149676 17040 149688
rect 17092 149676 17098 149728
rect 152734 149676 152740 149728
rect 152792 149716 152798 149728
rect 350534 149716 350540 149728
rect 152792 149688 350540 149716
rect 152792 149676 152798 149688
rect 350534 149676 350540 149688
rect 350592 149676 350598 149728
rect 6362 149064 6368 149116
rect 6420 149104 6426 149116
rect 8294 149104 8300 149116
rect 6420 149076 8300 149104
rect 6420 149064 6426 149076
rect 8294 149064 8300 149076
rect 8352 149064 8358 149116
rect 9122 149064 9128 149116
rect 9180 149104 9186 149116
rect 10226 149104 10232 149116
rect 9180 149076 10232 149104
rect 9180 149064 9186 149076
rect 10226 149064 10232 149076
rect 10284 149064 10290 149116
rect 14458 149064 14464 149116
rect 14516 149104 14522 149116
rect 15746 149104 15752 149116
rect 14516 149076 15752 149104
rect 14516 149064 14522 149076
rect 15746 149064 15752 149076
rect 15804 149064 15810 149116
rect 11974 147636 11980 147688
rect 12032 147676 12038 147688
rect 14274 147676 14280 147688
rect 12032 147648 14280 147676
rect 12032 147636 12038 147648
rect 14274 147636 14280 147648
rect 14332 147636 14338 147688
rect 151170 139340 151176 139392
rect 151228 139380 151234 139392
rect 580166 139380 580172 139392
rect 151228 139352 580172 139380
rect 151228 139340 151234 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 135804 3516 135856
rect 3568 135844 3574 135856
rect 4890 135844 4896 135856
rect 3568 135816 4896 135844
rect 3568 135804 3574 135816
rect 4890 135804 4896 135816
rect 4948 135804 4954 135856
rect 4890 134580 4896 134632
rect 4948 134620 4954 134632
rect 6178 134620 6184 134632
rect 4948 134592 6184 134620
rect 4948 134580 4954 134592
rect 6178 134580 6184 134592
rect 6236 134580 6242 134632
rect 156690 126896 156696 126948
rect 156748 126936 156754 126948
rect 580166 126936 580172 126948
rect 156748 126908 580172 126936
rect 156748 126896 156754 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 162118 113092 162124 113144
rect 162176 113132 162182 113144
rect 580166 113132 580172 113144
rect 162176 113104 580172 113132
rect 162176 113092 162182 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 151078 100648 151084 100700
rect 151136 100688 151142 100700
rect 580166 100688 580172 100700
rect 151136 100660 580172 100688
rect 151136 100648 151142 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3142 97928 3148 97980
rect 3200 97968 3206 97980
rect 18506 97968 18512 97980
rect 3200 97940 18512 97968
rect 3200 97928 3206 97940
rect 18506 97928 18512 97940
rect 18564 97928 18570 97980
rect 153930 86912 153936 86964
rect 153988 86952 153994 86964
rect 580166 86952 580172 86964
rect 153988 86924 580172 86952
rect 153988 86912 153994 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 2958 85484 2964 85536
rect 3016 85524 3022 85536
rect 12986 85524 12992 85536
rect 3016 85496 12992 85524
rect 3016 85484 3022 85496
rect 12986 85484 12992 85496
rect 13044 85484 13050 85536
rect 12986 82832 12992 82884
rect 13044 82872 13050 82884
rect 17126 82872 17132 82884
rect 13044 82844 17132 82872
rect 13044 82832 13050 82844
rect 17126 82832 17132 82844
rect 17184 82832 17190 82884
rect 152642 75828 152648 75880
rect 152700 75868 152706 75880
rect 156690 75868 156696 75880
rect 152700 75840 156696 75868
rect 152700 75828 152706 75840
rect 156690 75828 156696 75840
rect 156748 75828 156754 75880
rect 156598 74332 156604 74384
rect 156656 74372 156662 74384
rect 160094 74372 160100 74384
rect 156656 74344 160100 74372
rect 156656 74332 156662 74344
rect 160094 74332 160100 74344
rect 160152 74332 160158 74384
rect 160738 73108 160744 73160
rect 160796 73148 160802 73160
rect 579982 73148 579988 73160
rect 160796 73120 579988 73148
rect 160796 73108 160802 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 7558 71652 7564 71664
rect 3476 71624 7564 71652
rect 3476 71612 3482 71624
rect 7558 71612 7564 71624
rect 7616 71612 7622 71664
rect 576118 60664 576124 60716
rect 576176 60704 576182 60716
rect 580166 60704 580172 60716
rect 576176 60676 580172 60704
rect 576176 60664 576182 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3326 59304 3332 59356
rect 3384 59344 3390 59356
rect 10318 59344 10324 59356
rect 3384 59316 10324 59344
rect 3384 59304 3390 59316
rect 10318 59304 10324 59316
rect 10376 59304 10382 59356
rect 10318 56924 10324 56976
rect 10376 56964 10382 56976
rect 11698 56964 11704 56976
rect 10376 56936 11704 56964
rect 10376 56924 10382 56936
rect 11698 56924 11704 56936
rect 11756 56924 11762 56976
rect 152550 46860 152556 46912
rect 152608 46900 152614 46912
rect 580166 46900 580172 46912
rect 152608 46872 580172 46900
rect 152608 46860 152614 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 14366 45540 14372 45552
rect 3476 45512 14372 45540
rect 3476 45500 3482 45512
rect 14366 45500 14372 45512
rect 14424 45500 14430 45552
rect 278038 41012 278044 41064
rect 278096 41052 278102 41064
rect 282914 41052 282920 41064
rect 278096 41024 282920 41052
rect 278096 41012 278102 41024
rect 282914 41012 282920 41024
rect 282972 41012 282978 41064
rect 283558 39992 283564 40044
rect 283616 40032 283622 40044
rect 287790 40032 287796 40044
rect 283616 40004 287796 40032
rect 283616 39992 283622 40004
rect 287790 39992 287796 40004
rect 287848 39992 287854 40044
rect 287698 38564 287704 38616
rect 287756 38604 287762 38616
rect 295334 38604 295340 38616
rect 287756 38576 295340 38604
rect 287756 38564 287762 38576
rect 295334 38564 295340 38576
rect 295392 38564 295398 38616
rect 295978 36524 295984 36576
rect 296036 36564 296042 36576
rect 300670 36564 300676 36576
rect 296036 36536 300676 36564
rect 296036 36524 296042 36536
rect 300670 36524 300676 36536
rect 300728 36524 300734 36576
rect 282914 36252 282920 36304
rect 282972 36292 282978 36304
rect 287054 36292 287060 36304
rect 282972 36264 287060 36292
rect 282972 36252 282978 36264
rect 287054 36252 287060 36264
rect 287112 36252 287118 36304
rect 287790 35572 287796 35624
rect 287848 35612 287854 35624
rect 295426 35612 295432 35624
rect 287848 35584 295432 35612
rect 287848 35572 287854 35584
rect 295426 35572 295432 35584
rect 295484 35572 295490 35624
rect 300118 35028 300124 35080
rect 300176 35068 300182 35080
rect 303246 35068 303252 35080
rect 300176 35040 303252 35068
rect 300176 35028 300182 35040
rect 303246 35028 303252 35040
rect 303304 35028 303310 35080
rect 302878 33804 302884 33856
rect 302936 33844 302942 33856
rect 304994 33844 305000 33856
rect 302936 33816 305000 33844
rect 302936 33804 302942 33816
rect 304994 33804 305000 33816
rect 305052 33804 305058 33856
rect 295334 33736 295340 33788
rect 295392 33776 295398 33788
rect 299842 33776 299848 33788
rect 295392 33748 299848 33776
rect 295392 33736 295398 33748
rect 299842 33736 299848 33748
rect 299900 33736 299906 33788
rect 157978 33056 157984 33108
rect 158036 33096 158042 33108
rect 580166 33096 580172 33108
rect 158036 33068 580172 33096
rect 158036 33056 158042 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 32580 3424 32632
rect 3476 32620 3482 32632
rect 8938 32620 8944 32632
rect 3476 32592 8944 32620
rect 3476 32580 3482 32592
rect 8938 32580 8944 32592
rect 8996 32580 9002 32632
rect 300670 32580 300676 32632
rect 300728 32620 300734 32632
rect 302510 32620 302516 32632
rect 300728 32592 302516 32620
rect 300728 32580 300734 32592
rect 302510 32580 302516 32592
rect 302568 32580 302574 32632
rect 152458 32376 152464 32428
rect 152516 32416 152522 32428
rect 165890 32416 165896 32428
rect 152516 32388 165896 32416
rect 152516 32376 152522 32388
rect 165890 32376 165896 32388
rect 165948 32376 165954 32428
rect 305638 32376 305644 32428
rect 305696 32416 305702 32428
rect 309226 32416 309232 32428
rect 305696 32388 309232 32416
rect 305696 32376 305702 32388
rect 309226 32376 309232 32388
rect 309284 32376 309290 32428
rect 287054 31696 287060 31748
rect 287112 31736 287118 31748
rect 295334 31736 295340 31748
rect 287112 31708 295340 31736
rect 287112 31696 287118 31708
rect 295334 31696 295340 31708
rect 295392 31696 295398 31748
rect 303246 31696 303252 31748
rect 303304 31736 303310 31748
rect 305086 31736 305092 31748
rect 303304 31708 305092 31736
rect 303304 31696 303310 31708
rect 305086 31696 305092 31708
rect 305144 31696 305150 31748
rect 166258 31356 166264 31408
rect 166316 31396 166322 31408
rect 168466 31396 168472 31408
rect 166316 31368 168472 31396
rect 166316 31356 166322 31368
rect 168466 31356 168472 31368
rect 168524 31356 168530 31408
rect 153838 31084 153844 31136
rect 153896 31124 153902 31136
rect 179414 31124 179420 31136
rect 153896 31096 179420 31124
rect 153896 31084 153902 31096
rect 179414 31084 179420 31096
rect 179472 31084 179478 31136
rect 156690 31016 156696 31068
rect 156748 31056 156754 31068
rect 216030 31056 216036 31068
rect 156748 31028 216036 31056
rect 156748 31016 156754 31028
rect 216030 31016 216036 31028
rect 216088 31016 216094 31068
rect 309778 31016 309784 31068
rect 309836 31056 309842 31068
rect 328086 31056 328092 31068
rect 309836 31028 328092 31056
rect 309836 31016 309842 31028
rect 328086 31016 328092 31028
rect 328144 31016 328150 31068
rect 165890 30268 165896 30320
rect 165948 30308 165954 30320
rect 172514 30308 172520 30320
rect 165948 30280 172520 30308
rect 165948 30268 165954 30280
rect 172514 30268 172520 30280
rect 172572 30268 172578 30320
rect 215938 30268 215944 30320
rect 215996 30308 216002 30320
rect 218054 30308 218060 30320
rect 215996 30280 218060 30308
rect 215996 30268 216002 30280
rect 218054 30268 218060 30280
rect 218112 30268 218118 30320
rect 233878 30268 233884 30320
rect 233936 30308 233942 30320
rect 235994 30308 236000 30320
rect 233936 30280 236000 30308
rect 233936 30268 233942 30280
rect 235994 30268 236000 30280
rect 236052 30268 236058 30320
rect 238018 30268 238024 30320
rect 238076 30308 238082 30320
rect 240134 30308 240140 30320
rect 238076 30280 240140 30308
rect 238076 30268 238082 30280
rect 240134 30268 240140 30280
rect 240192 30268 240198 30320
rect 385678 30268 385684 30320
rect 385736 30308 385742 30320
rect 388530 30308 388536 30320
rect 385736 30280 388536 30308
rect 385736 30268 385742 30280
rect 388530 30268 388536 30280
rect 388588 30268 388594 30320
rect 327718 29724 327724 29776
rect 327776 29764 327782 29776
rect 341610 29764 341616 29776
rect 327776 29736 341616 29764
rect 327776 29724 327782 29736
rect 341610 29724 341616 29736
rect 341668 29724 341674 29776
rect 304994 29656 305000 29708
rect 305052 29696 305058 29708
rect 327810 29696 327816 29708
rect 305052 29668 327816 29696
rect 305052 29656 305058 29668
rect 327810 29656 327816 29668
rect 327868 29656 327874 29708
rect 180058 29588 180064 29640
rect 180116 29628 180122 29640
rect 193306 29628 193312 29640
rect 180116 29600 193312 29628
rect 180116 29588 180122 29600
rect 193306 29588 193312 29600
rect 193364 29588 193370 29640
rect 246298 29588 246304 29640
rect 246356 29628 246362 29640
rect 253934 29628 253940 29640
rect 246356 29600 253940 29628
rect 246356 29588 246362 29600
rect 253934 29588 253940 29600
rect 253992 29588 253998 29640
rect 295426 29588 295432 29640
rect 295484 29628 295490 29640
rect 354030 29628 354036 29640
rect 295484 29600 354036 29628
rect 295484 29588 295490 29600
rect 354030 29588 354036 29600
rect 354088 29588 354094 29640
rect 220078 28908 220084 28960
rect 220136 28948 220142 28960
rect 222194 28948 222200 28960
rect 220136 28920 222200 28948
rect 220136 28908 220142 28920
rect 222194 28908 222200 28920
rect 222252 28908 222258 28960
rect 328086 28568 328092 28620
rect 328144 28608 328150 28620
rect 336090 28608 336096 28620
rect 328144 28580 336096 28608
rect 328144 28568 328150 28580
rect 336090 28568 336096 28580
rect 336148 28568 336154 28620
rect 299842 28500 299848 28552
rect 299900 28540 299906 28552
rect 349798 28540 349804 28552
rect 299900 28512 349804 28540
rect 299900 28500 299906 28512
rect 349798 28500 349804 28512
rect 349856 28500 349862 28552
rect 353938 28500 353944 28552
rect 353996 28540 354002 28552
rect 381630 28540 381636 28552
rect 353996 28512 381636 28540
rect 353996 28500 354002 28512
rect 381630 28500 381636 28512
rect 381688 28500 381694 28552
rect 305086 28432 305092 28484
rect 305144 28472 305150 28484
rect 359550 28472 359556 28484
rect 305144 28444 359556 28472
rect 305144 28432 305150 28444
rect 359550 28432 359556 28444
rect 359608 28432 359614 28484
rect 302510 28364 302516 28416
rect 302568 28404 302574 28416
rect 377950 28404 377956 28416
rect 302568 28376 377956 28404
rect 302568 28364 302574 28376
rect 377950 28364 377956 28376
rect 378008 28364 378014 28416
rect 295334 28296 295340 28348
rect 295392 28336 295398 28348
rect 371878 28336 371884 28348
rect 295392 28308 371884 28336
rect 295392 28296 295398 28308
rect 371878 28296 371884 28308
rect 371936 28296 371942 28348
rect 388438 28296 388444 28348
rect 388496 28336 388502 28348
rect 400030 28336 400036 28348
rect 388496 28308 400036 28336
rect 388496 28296 388502 28308
rect 400030 28296 400036 28308
rect 400088 28296 400094 28348
rect 309226 28228 309232 28280
rect 309284 28268 309290 28280
rect 395338 28268 395344 28280
rect 309284 28240 395344 28268
rect 309284 28228 309290 28240
rect 395338 28228 395344 28240
rect 395396 28228 395402 28280
rect 406378 27548 406384 27600
rect 406436 27588 406442 27600
rect 409046 27588 409052 27600
rect 406436 27560 409052 27588
rect 406436 27548 406442 27560
rect 409046 27548 409052 27560
rect 409104 27548 409110 27600
rect 17034 27072 17040 27124
rect 17092 27112 17098 27124
rect 17310 27112 17316 27124
rect 17092 27084 17316 27112
rect 17092 27072 17098 27084
rect 17310 27072 17316 27084
rect 17368 27072 17374 27124
rect 17494 26732 17500 26784
rect 17552 26772 17558 26784
rect 17678 26772 17684 26784
rect 17552 26744 17684 26772
rect 17552 26732 17558 26744
rect 17678 26732 17684 26744
rect 17736 26732 17742 26784
rect 153286 26664 153292 26716
rect 153344 26704 153350 26716
rect 255958 26704 255964 26716
rect 153344 26676 255964 26704
rect 153344 26664 153350 26676
rect 255958 26664 255964 26676
rect 256016 26664 256022 26716
rect 157242 26596 157248 26648
rect 157300 26636 157306 26648
rect 291838 26636 291844 26648
rect 157300 26608 291844 26636
rect 157300 26596 157306 26608
rect 291838 26596 291844 26608
rect 291896 26596 291902 26648
rect 152090 26528 152096 26580
rect 152148 26568 152154 26580
rect 318058 26568 318064 26580
rect 152148 26540 318064 26568
rect 152148 26528 152154 26540
rect 318058 26528 318064 26540
rect 318116 26528 318122 26580
rect 159358 26460 159364 26512
rect 159416 26500 159422 26512
rect 345014 26500 345020 26512
rect 159416 26472 345020 26500
rect 159416 26460 159422 26472
rect 345014 26460 345020 26472
rect 345072 26460 345078 26512
rect 157334 26392 157340 26444
rect 157392 26432 157398 26444
rect 355318 26432 355324 26444
rect 157392 26404 355324 26432
rect 157392 26392 157398 26404
rect 355318 26392 355324 26404
rect 355376 26392 355382 26444
rect 156966 26324 156972 26376
rect 157024 26364 157030 26376
rect 509878 26364 509884 26376
rect 157024 26336 509884 26364
rect 157024 26324 157030 26336
rect 509878 26324 509884 26336
rect 509936 26324 509942 26376
rect 154942 26256 154948 26308
rect 155000 26296 155006 26308
rect 510614 26296 510620 26308
rect 155000 26268 510620 26296
rect 155000 26256 155006 26268
rect 510614 26256 510620 26268
rect 510672 26256 510678 26308
rect 409138 26052 409144 26104
rect 409196 26092 409202 26104
rect 413462 26092 413468 26104
rect 409196 26064 413468 26092
rect 409196 26052 409202 26064
rect 413462 26052 413468 26064
rect 413520 26052 413526 26104
rect 341610 25916 341616 25968
rect 341668 25956 341674 25968
rect 346302 25956 346308 25968
rect 341668 25928 346308 25956
rect 341668 25916 341674 25928
rect 346302 25916 346308 25928
rect 346360 25916 346366 25968
rect 371878 25576 371884 25628
rect 371936 25616 371942 25628
rect 380894 25616 380900 25628
rect 371936 25588 380900 25616
rect 371936 25576 371942 25588
rect 380894 25576 380900 25588
rect 380952 25576 380958 25628
rect 345014 25508 345020 25560
rect 345072 25548 345078 25560
rect 485038 25548 485044 25560
rect 345072 25520 485044 25548
rect 345072 25508 345078 25520
rect 485038 25508 485044 25520
rect 485096 25508 485102 25560
rect 160186 25304 160192 25356
rect 160244 25344 160250 25356
rect 303614 25344 303620 25356
rect 160244 25316 303620 25344
rect 160244 25304 160250 25316
rect 303614 25304 303620 25316
rect 303672 25304 303678 25356
rect 153378 25236 153384 25288
rect 153436 25276 153442 25288
rect 327994 25276 328000 25288
rect 153436 25248 328000 25276
rect 153436 25236 153442 25248
rect 327994 25236 328000 25248
rect 328052 25236 328058 25288
rect 156046 25168 156052 25220
rect 156104 25208 156110 25220
rect 355870 25208 355876 25220
rect 156104 25180 355876 25208
rect 156104 25168 156110 25180
rect 355870 25168 355876 25180
rect 355928 25168 355934 25220
rect 156598 25100 156604 25152
rect 156656 25140 156662 25152
rect 403894 25140 403900 25152
rect 156656 25112 403900 25140
rect 156656 25100 156662 25112
rect 403894 25100 403900 25112
rect 403952 25100 403958 25152
rect 152918 25032 152924 25084
rect 152976 25072 152982 25084
rect 445754 25072 445760 25084
rect 152976 25044 445760 25072
rect 152976 25032 152982 25044
rect 445754 25032 445760 25044
rect 445812 25032 445818 25084
rect 157886 24964 157892 25016
rect 157944 25004 157950 25016
rect 488534 25004 488540 25016
rect 157944 24976 488540 25004
rect 157944 24964 157950 24976
rect 488534 24964 488540 24976
rect 488592 24964 488598 25016
rect 159450 24896 159456 24948
rect 159508 24936 159514 24948
rect 494698 24936 494704 24948
rect 159508 24908 494704 24936
rect 159508 24896 159514 24908
rect 494698 24896 494704 24908
rect 494756 24896 494762 24948
rect 153102 24828 153108 24880
rect 153160 24868 153166 24880
rect 556154 24868 556160 24880
rect 153160 24840 556160 24868
rect 153160 24828 153166 24840
rect 556154 24828 556160 24840
rect 556212 24828 556218 24880
rect 388530 24624 388536 24676
rect 388588 24664 388594 24676
rect 391290 24664 391296 24676
rect 388588 24636 391296 24664
rect 388588 24624 388594 24636
rect 391290 24624 391296 24636
rect 391348 24624 391354 24676
rect 188338 24148 188344 24200
rect 188396 24188 188402 24200
rect 190454 24188 190460 24200
rect 188396 24160 190460 24188
rect 188396 24148 188402 24160
rect 190454 24148 190460 24160
rect 190512 24148 190518 24200
rect 381538 24148 381544 24200
rect 381596 24188 381602 24200
rect 388346 24188 388352 24200
rect 381596 24160 388352 24188
rect 381596 24148 381602 24160
rect 388346 24148 388352 24160
rect 388404 24148 388410 24200
rect 303614 24080 303620 24132
rect 303672 24120 303678 24132
rect 549254 24120 549260 24132
rect 303672 24092 549260 24120
rect 303672 24080 303678 24092
rect 549254 24080 549260 24092
rect 549312 24080 549318 24132
rect 159542 23944 159548 23996
rect 159600 23984 159606 23996
rect 215294 23984 215300 23996
rect 159600 23956 215300 23984
rect 159600 23944 159606 23956
rect 215294 23944 215300 23956
rect 215352 23944 215358 23996
rect 158070 23876 158076 23928
rect 158128 23916 158134 23928
rect 254026 23916 254032 23928
rect 158128 23888 254032 23916
rect 158128 23876 158134 23888
rect 254026 23876 254032 23888
rect 254084 23876 254090 23928
rect 155770 23808 155776 23860
rect 155828 23848 155834 23860
rect 305638 23848 305644 23860
rect 155828 23820 305644 23848
rect 155828 23808 155834 23820
rect 305638 23808 305644 23820
rect 305696 23808 305702 23860
rect 152826 23740 152832 23792
rect 152884 23780 152890 23792
rect 309134 23780 309140 23792
rect 152884 23752 309140 23780
rect 152884 23740 152890 23752
rect 309134 23740 309140 23752
rect 309192 23740 309198 23792
rect 403618 23740 403624 23792
rect 403676 23780 403682 23792
rect 406654 23780 406660 23792
rect 403676 23752 406660 23780
rect 403676 23740 403682 23752
rect 406654 23740 406660 23752
rect 406712 23740 406718 23792
rect 553394 23712 553400 23724
rect 153212 23684 553400 23712
rect 152642 23400 152648 23452
rect 152700 23440 152706 23452
rect 153212 23440 153240 23684
rect 553394 23672 553400 23684
rect 553452 23672 553458 23724
rect 156690 23604 156696 23656
rect 156748 23644 156754 23656
rect 563054 23644 563060 23656
rect 156748 23616 563060 23644
rect 156748 23604 156754 23616
rect 563054 23604 563060 23616
rect 563112 23604 563118 23656
rect 157058 23536 157064 23588
rect 157116 23576 157122 23588
rect 571334 23576 571340 23588
rect 157116 23548 571340 23576
rect 157116 23536 157122 23548
rect 571334 23536 571340 23548
rect 571392 23536 571398 23588
rect 155126 23468 155132 23520
rect 155184 23508 155190 23520
rect 575474 23508 575480 23520
rect 155184 23480 575480 23508
rect 155184 23468 155190 23480
rect 575474 23468 575480 23480
rect 575532 23468 575538 23520
rect 152700 23412 153240 23440
rect 152700 23400 152706 23412
rect 341518 23400 341524 23452
rect 341576 23440 341582 23452
rect 345750 23440 345756 23452
rect 341576 23412 345756 23440
rect 341576 23400 341582 23412
rect 345750 23400 345756 23412
rect 345808 23400 345814 23452
rect 399478 23400 399484 23452
rect 399536 23440 399542 23452
rect 403618 23440 403624 23452
rect 399536 23412 403624 23440
rect 399536 23400 399542 23412
rect 403618 23400 403624 23412
rect 403676 23400 403682 23452
rect 462958 23400 462964 23452
rect 463016 23440 463022 23452
rect 466730 23440 466736 23452
rect 463016 23412 466736 23440
rect 463016 23400 463022 23412
rect 466730 23400 466736 23412
rect 466788 23400 466794 23452
rect 335998 23264 336004 23316
rect 336056 23304 336062 23316
rect 341610 23304 341616 23316
rect 336056 23276 341616 23304
rect 336056 23264 336062 23276
rect 341610 23264 341616 23276
rect 341668 23264 341674 23316
rect 453298 23128 453304 23180
rect 453356 23168 453362 23180
rect 458174 23168 458180 23180
rect 453356 23140 458180 23168
rect 453356 23128 453362 23140
rect 458174 23128 458180 23140
rect 458232 23128 458238 23180
rect 359458 22992 359464 23044
rect 359516 23032 359522 23044
rect 363690 23032 363696 23044
rect 359516 23004 363696 23032
rect 359516 22992 359522 23004
rect 363690 22992 363696 23004
rect 363748 22992 363754 23044
rect 409046 22992 409052 23044
rect 409104 23032 409110 23044
rect 417510 23032 417516 23044
rect 409104 23004 417516 23032
rect 409104 22992 409110 23004
rect 417510 22992 417516 23004
rect 417568 22992 417574 23044
rect 421558 22992 421564 23044
rect 421616 23032 421622 23044
rect 426802 23032 426808 23044
rect 421616 23004 426808 23032
rect 421616 22992 421622 23004
rect 426802 22992 426808 23004
rect 426860 22992 426866 23044
rect 345658 22924 345664 22976
rect 345716 22964 345722 22976
rect 356790 22964 356796 22976
rect 345716 22936 356796 22964
rect 345716 22924 345722 22936
rect 356790 22924 356796 22936
rect 356848 22924 356854 22976
rect 371970 22924 371976 22976
rect 372028 22964 372034 22976
rect 378042 22964 378048 22976
rect 372028 22936 378048 22964
rect 372028 22924 372034 22936
rect 378042 22924 378048 22936
rect 378100 22924 378106 22976
rect 150894 22856 150900 22908
rect 150952 22896 150958 22908
rect 152090 22896 152096 22908
rect 150952 22868 152096 22896
rect 150952 22856 150958 22868
rect 152090 22856 152096 22868
rect 152148 22856 152154 22908
rect 255958 22856 255964 22908
rect 256016 22896 256022 22908
rect 334618 22896 334624 22908
rect 256016 22868 334624 22896
rect 256016 22856 256022 22868
rect 334618 22856 334624 22868
rect 334676 22856 334682 22908
rect 346302 22856 346308 22908
rect 346360 22896 346366 22908
rect 371234 22896 371240 22908
rect 346360 22868 371240 22896
rect 346360 22856 346366 22868
rect 371234 22856 371240 22868
rect 371292 22856 371298 22908
rect 377950 22856 377956 22908
rect 378008 22896 378014 22908
rect 388530 22896 388536 22908
rect 378008 22868 388536 22896
rect 378008 22856 378014 22868
rect 388530 22856 388536 22868
rect 388588 22856 388594 22908
rect 391198 22856 391204 22908
rect 391256 22896 391262 22908
rect 408586 22896 408592 22908
rect 391256 22868 408592 22896
rect 391256 22856 391262 22868
rect 408586 22856 408592 22868
rect 408644 22856 408650 22908
rect 417418 22856 417424 22908
rect 417476 22896 417482 22908
rect 430574 22896 430580 22908
rect 417476 22868 430580 22896
rect 417476 22856 417482 22868
rect 430574 22856 430580 22868
rect 430632 22856 430638 22908
rect 216030 22788 216036 22840
rect 216088 22828 216094 22840
rect 218146 22828 218152 22840
rect 216088 22800 218152 22828
rect 216088 22788 216094 22800
rect 218146 22788 218152 22800
rect 218204 22788 218210 22840
rect 327994 22788 328000 22840
rect 328052 22828 328058 22840
rect 480898 22828 480904 22840
rect 328052 22800 480904 22828
rect 328052 22788 328058 22800
rect 480898 22788 480904 22800
rect 480956 22788 480962 22840
rect 215294 22720 215300 22772
rect 215352 22760 215358 22772
rect 471422 22760 471428 22772
rect 215352 22732 471428 22760
rect 215352 22720 215358 22732
rect 471422 22720 471428 22732
rect 471480 22720 471486 22772
rect 151354 22652 151360 22704
rect 151412 22692 151418 22704
rect 176746 22692 176752 22704
rect 151412 22664 176752 22692
rect 151412 22652 151418 22664
rect 176746 22652 176752 22664
rect 176804 22652 176810 22704
rect 157426 22584 157432 22636
rect 157484 22624 157490 22636
rect 241422 22624 241428 22636
rect 157484 22596 241428 22624
rect 157484 22584 157490 22596
rect 241422 22584 241428 22596
rect 241480 22584 241486 22636
rect 154022 22516 154028 22568
rect 154080 22556 154086 22568
rect 284294 22556 284300 22568
rect 154080 22528 284300 22556
rect 154080 22516 154086 22528
rect 284294 22516 284300 22528
rect 284352 22516 284358 22568
rect 154206 22448 154212 22500
rect 154264 22488 154270 22500
rect 327074 22488 327080 22500
rect 154264 22460 327080 22488
rect 154264 22448 154270 22460
rect 327074 22448 327080 22460
rect 327132 22448 327138 22500
rect 153010 22380 153016 22432
rect 153068 22420 153074 22432
rect 345842 22420 345848 22432
rect 153068 22392 345848 22420
rect 153068 22380 153074 22392
rect 345842 22380 345848 22392
rect 345900 22380 345906 22432
rect 156506 22312 156512 22364
rect 156564 22352 156570 22364
rect 399570 22352 399576 22364
rect 156564 22324 399576 22352
rect 156564 22312 156570 22324
rect 399570 22312 399576 22324
rect 399628 22312 399634 22364
rect 413462 22312 413468 22364
rect 413520 22352 413526 22364
rect 421006 22352 421012 22364
rect 413520 22324 421012 22352
rect 413520 22312 413526 22324
rect 421006 22312 421012 22324
rect 421064 22312 421070 22364
rect 154298 22244 154304 22296
rect 154356 22284 154362 22296
rect 438854 22284 438860 22296
rect 154356 22256 438860 22284
rect 154356 22244 154362 22256
rect 438854 22244 438860 22256
rect 438912 22244 438918 22296
rect 153930 22176 153936 22228
rect 153988 22216 153994 22228
rect 567194 22216 567200 22228
rect 153988 22188 567200 22216
rect 153988 22176 153994 22188
rect 567194 22176 567200 22188
rect 567252 22176 567258 22228
rect 150986 22108 150992 22160
rect 151044 22148 151050 22160
rect 153102 22148 153108 22160
rect 151044 22120 153108 22148
rect 151044 22108 151050 22120
rect 153102 22108 153108 22120
rect 153160 22108 153166 22160
rect 158162 22108 158168 22160
rect 158220 22148 158226 22160
rect 574094 22148 574100 22160
rect 158220 22120 574100 22148
rect 158220 22108 158226 22120
rect 574094 22108 574100 22120
rect 574152 22108 574158 22160
rect 241422 21428 241428 21480
rect 241480 21468 241486 21480
rect 288434 21468 288440 21480
rect 241480 21440 288440 21468
rect 241480 21428 241486 21440
rect 288434 21428 288440 21440
rect 288492 21428 288498 21480
rect 355870 21428 355876 21480
rect 355928 21468 355934 21480
rect 370498 21468 370504 21480
rect 355928 21440 370504 21468
rect 355928 21428 355934 21440
rect 370498 21428 370504 21440
rect 370556 21428 370562 21480
rect 155954 21360 155960 21412
rect 156012 21400 156018 21412
rect 157886 21400 157892 21412
rect 156012 21372 157892 21400
rect 156012 21360 156018 21372
rect 157886 21360 157892 21372
rect 157944 21360 157950 21412
rect 284294 21360 284300 21412
rect 284352 21400 284358 21412
rect 424962 21400 424968 21412
rect 284352 21372 424968 21400
rect 284352 21360 284358 21372
rect 424962 21360 424968 21372
rect 425020 21360 425026 21412
rect 155678 21292 155684 21344
rect 155736 21332 155742 21344
rect 157058 21332 157064 21344
rect 155736 21304 157064 21332
rect 155736 21292 155742 21304
rect 157058 21292 157064 21304
rect 157116 21292 157122 21344
rect 158254 21292 158260 21344
rect 158312 21332 158318 21344
rect 160186 21332 160192 21344
rect 158312 21304 160192 21332
rect 158312 21292 158318 21304
rect 160186 21292 160192 21304
rect 160244 21292 160250 21344
rect 153838 21224 153844 21276
rect 153896 21264 153902 21276
rect 215294 21264 215300 21276
rect 153896 21236 215300 21264
rect 153896 21224 153902 21236
rect 215294 21224 215300 21236
rect 215352 21224 215358 21276
rect 154390 21156 154396 21208
rect 154448 21196 154454 21208
rect 241422 21196 241428 21208
rect 154448 21168 241428 21196
rect 154448 21156 154454 21168
rect 241422 21156 241428 21168
rect 241480 21156 241486 21208
rect 155862 21088 155868 21140
rect 155920 21128 155926 21140
rect 260742 21128 260748 21140
rect 155920 21100 260748 21128
rect 155920 21088 155926 21100
rect 260742 21088 260748 21100
rect 260800 21088 260806 21140
rect 151446 21020 151452 21072
rect 151504 21060 151510 21072
rect 300762 21060 300768 21072
rect 151504 21032 300768 21060
rect 151504 21020 151510 21032
rect 300762 21020 300768 21032
rect 300820 21020 300826 21072
rect 152550 20952 152556 21004
rect 152608 20992 152614 21004
rect 319530 20992 319536 21004
rect 152608 20964 319536 20992
rect 152608 20952 152614 20964
rect 319530 20952 319536 20964
rect 319588 20952 319594 21004
rect 151998 20884 152004 20936
rect 152056 20924 152062 20936
rect 155126 20924 155132 20936
rect 152056 20896 155132 20924
rect 152056 20884 152062 20896
rect 155126 20884 155132 20896
rect 155184 20884 155190 20936
rect 155218 20884 155224 20936
rect 155276 20924 155282 20936
rect 157242 20924 157248 20936
rect 155276 20896 157248 20924
rect 155276 20884 155282 20896
rect 157242 20884 157248 20896
rect 157300 20884 157306 20936
rect 413922 20924 413928 20936
rect 157352 20896 413928 20924
rect 154482 20816 154488 20868
rect 154540 20856 154546 20868
rect 157352 20856 157380 20896
rect 413922 20884 413928 20896
rect 413980 20884 413986 20936
rect 507118 20856 507124 20868
rect 154540 20828 157380 20856
rect 157444 20828 507124 20856
rect 154540 20816 154546 20828
rect 154114 20748 154120 20800
rect 154172 20788 154178 20800
rect 157444 20788 157472 20828
rect 507118 20816 507124 20828
rect 507176 20816 507182 20868
rect 534718 20788 534724 20800
rect 154172 20760 157472 20788
rect 157536 20760 534724 20788
rect 154172 20748 154178 20760
rect 153286 20720 153292 20732
rect 151786 20692 153292 20720
rect 15930 20612 15936 20664
rect 15988 20652 15994 20664
rect 18506 20652 18512 20664
rect 15988 20624 18512 20652
rect 15988 20612 15994 20624
rect 18506 20612 18512 20624
rect 18564 20612 18570 20664
rect 19058 20612 19064 20664
rect 19116 20652 19122 20664
rect 19794 20652 19800 20664
rect 19116 20624 19800 20652
rect 19116 20612 19122 20624
rect 19794 20612 19800 20624
rect 19852 20612 19858 20664
rect 151262 20612 151268 20664
rect 151320 20652 151326 20664
rect 151786 20652 151814 20692
rect 153286 20680 153292 20692
rect 153344 20680 153350 20732
rect 157536 20720 157564 20760
rect 534718 20748 534724 20760
rect 534776 20748 534782 20800
rect 154592 20692 157564 20720
rect 151320 20624 151814 20652
rect 151320 20612 151326 20624
rect 152366 20612 152372 20664
rect 152424 20652 152430 20664
rect 154592 20652 154620 20692
rect 157978 20680 157984 20732
rect 158036 20720 158042 20732
rect 552014 20720 552020 20732
rect 158036 20692 552020 20720
rect 158036 20680 158042 20692
rect 552014 20680 552020 20692
rect 552072 20680 552078 20732
rect 152424 20624 154620 20652
rect 152424 20612 152430 20624
rect 406654 20612 406660 20664
rect 406712 20652 406718 20664
rect 413278 20652 413284 20664
rect 406712 20624 413284 20652
rect 406712 20612 406718 20624
rect 413278 20612 413284 20624
rect 413336 20612 413342 20664
rect 466730 20612 466736 20664
rect 466788 20652 466794 20664
rect 471330 20652 471336 20664
rect 466788 20624 471336 20652
rect 466788 20612 466794 20624
rect 471330 20612 471336 20624
rect 471388 20612 471394 20664
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 17678 20584 17684 20596
rect 13136 20556 17684 20584
rect 13136 20544 13142 20556
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 153286 20544 153292 20596
rect 153344 20584 153350 20596
rect 154942 20584 154948 20596
rect 153344 20556 154948 20584
rect 153344 20544 153350 20556
rect 154942 20544 154948 20556
rect 155000 20544 155006 20596
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 17126 20516 17132 20528
rect 13044 20488 17132 20516
rect 13044 20476 13050 20488
rect 17126 20476 17132 20488
rect 17184 20476 17190 20528
rect 151538 20272 151544 20324
rect 151596 20312 151602 20324
rect 152918 20312 152924 20324
rect 151596 20284 152924 20312
rect 151596 20272 151602 20284
rect 152918 20272 152924 20284
rect 152976 20272 152982 20324
rect 155494 20136 155500 20188
rect 155552 20176 155558 20188
rect 156966 20176 156972 20188
rect 155552 20148 156972 20176
rect 155552 20136 155558 20148
rect 156966 20136 156972 20148
rect 157024 20136 157030 20188
rect 380894 20136 380900 20188
rect 380952 20176 380958 20188
rect 399478 20176 399484 20188
rect 380952 20148 399484 20176
rect 380952 20136 380958 20148
rect 399478 20136 399484 20148
rect 399536 20136 399542 20188
rect 400030 20136 400036 20188
rect 400088 20176 400094 20188
rect 407022 20176 407028 20188
rect 400088 20148 407028 20176
rect 400088 20136 400094 20148
rect 407022 20136 407028 20148
rect 407080 20136 407086 20188
rect 430574 20136 430580 20188
rect 430632 20176 430638 20188
rect 435542 20176 435548 20188
rect 430632 20148 435548 20176
rect 430632 20136 430638 20148
rect 435542 20136 435548 20148
rect 435600 20136 435606 20188
rect 439498 20136 439504 20188
rect 439556 20176 439562 20188
rect 453298 20176 453304 20188
rect 439556 20148 453304 20176
rect 439556 20136 439562 20148
rect 453298 20136 453304 20148
rect 453356 20136 453362 20188
rect 458174 20136 458180 20188
rect 458232 20176 458238 20188
rect 467190 20176 467196 20188
rect 458232 20148 467196 20176
rect 458232 20136 458238 20148
rect 467190 20136 467196 20148
rect 467248 20136 467254 20188
rect 13262 20068 13268 20120
rect 13320 20108 13326 20120
rect 19702 20108 19708 20120
rect 13320 20080 19708 20108
rect 13320 20068 13326 20080
rect 19702 20068 19708 20080
rect 19760 20068 19766 20120
rect 153102 20068 153108 20120
rect 153160 20108 153166 20120
rect 156598 20108 156604 20120
rect 153160 20080 156604 20108
rect 153160 20068 153166 20080
rect 156598 20068 156604 20080
rect 156656 20068 156662 20120
rect 327810 20068 327816 20120
rect 327868 20108 327874 20120
rect 335998 20108 336004 20120
rect 327868 20080 336004 20108
rect 327868 20068 327874 20080
rect 335998 20068 336004 20080
rect 336056 20068 336062 20120
rect 371234 20068 371240 20120
rect 371292 20108 371298 20120
rect 377582 20108 377588 20120
rect 371292 20080 377588 20108
rect 371292 20068 371298 20080
rect 377582 20068 377588 20080
rect 377640 20068 377646 20120
rect 378042 20068 378048 20120
rect 378100 20108 378106 20120
rect 403710 20108 403716 20120
rect 378100 20080 403716 20108
rect 378100 20068 378106 20080
rect 403710 20068 403716 20080
rect 403768 20068 403774 20120
rect 413922 20068 413928 20120
rect 413980 20108 413986 20120
rect 495434 20108 495440 20120
rect 413980 20080 495440 20108
rect 413980 20068 413986 20080
rect 495434 20068 495440 20080
rect 495492 20068 495498 20120
rect 3142 20000 3148 20052
rect 3200 20040 3206 20052
rect 4798 20040 4804 20052
rect 3200 20012 4804 20040
rect 3200 20000 3206 20012
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 19610 20040 19616 20052
rect 11940 20012 19616 20040
rect 11940 20000 11946 20012
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 152734 20000 152740 20052
rect 152792 20040 152798 20052
rect 157794 20040 157800 20052
rect 152792 20012 157800 20040
rect 152792 20000 152798 20012
rect 157794 20000 157800 20012
rect 157852 20000 157858 20052
rect 300762 20000 300768 20052
rect 300820 20040 300826 20052
rect 499574 20040 499580 20052
rect 300820 20012 499580 20040
rect 300820 20000 300826 20012
rect 499574 20000 499580 20012
rect 499632 20000 499638 20052
rect 6362 19932 6368 19984
rect 6420 19972 6426 19984
rect 19886 19972 19892 19984
rect 6420 19944 19892 19972
rect 6420 19932 6426 19944
rect 19886 19932 19892 19944
rect 19944 19932 19950 19984
rect 151078 19932 151084 19984
rect 151136 19972 151142 19984
rect 155862 19972 155868 19984
rect 151136 19944 155868 19972
rect 151136 19932 151142 19944
rect 155862 19932 155868 19944
rect 155920 19932 155926 19984
rect 215294 19932 215300 19984
rect 215352 19972 215358 19984
rect 222930 19972 222936 19984
rect 215352 19944 222936 19972
rect 215352 19932 215358 19944
rect 222930 19932 222936 19944
rect 222988 19932 222994 19984
rect 241422 19932 241428 19984
rect 241480 19972 241486 19984
rect 542354 19972 542360 19984
rect 241480 19944 542360 19972
rect 241480 19932 241486 19944
rect 542354 19932 542360 19944
rect 542412 19932 542418 19984
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 3660 19876 66484 19904
rect 3660 19864 3666 19876
rect 66456 19848 66484 19876
rect 84166 19876 103514 19904
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 17828 19808 60734 19836
rect 17828 19796 17834 19808
rect 10410 19728 10416 19780
rect 10468 19768 10474 19780
rect 35802 19768 35808 19780
rect 10468 19740 35808 19768
rect 10468 19728 10474 19740
rect 35802 19728 35808 19740
rect 35860 19728 35866 19780
rect 17034 19660 17040 19712
rect 17092 19700 17098 19712
rect 23474 19700 23480 19712
rect 17092 19672 23480 19700
rect 17092 19660 17098 19672
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 60706 19700 60734 19808
rect 66438 19796 66444 19848
rect 66496 19796 66502 19848
rect 70670 19700 70676 19712
rect 60706 19672 70676 19700
rect 70670 19660 70676 19672
rect 70728 19660 70734 19712
rect 81434 19660 81440 19712
rect 81492 19700 81498 19712
rect 84166 19700 84194 19876
rect 95234 19796 95240 19848
rect 95292 19836 95298 19848
rect 95924 19836 95930 19848
rect 95292 19808 95930 19836
rect 95292 19796 95298 19808
rect 95924 19796 95930 19808
rect 95982 19796 95988 19848
rect 100938 19796 100944 19848
rect 100996 19836 101002 19848
rect 101996 19836 102002 19848
rect 100996 19808 102002 19836
rect 100996 19796 101002 19808
rect 101996 19796 102002 19808
rect 102054 19796 102060 19848
rect 81492 19672 84194 19700
rect 103486 19700 103514 19876
rect 119844 19864 119850 19916
rect 119902 19904 119908 19916
rect 150894 19904 150900 19916
rect 119902 19876 122834 19904
rect 119902 19864 119908 19876
rect 109218 19796 109224 19848
rect 109276 19836 109282 19848
rect 110276 19836 110282 19848
rect 109276 19808 110282 19836
rect 109276 19796 109282 19808
rect 110276 19796 110282 19808
rect 110334 19796 110340 19848
rect 111978 19796 111984 19848
rect 112036 19836 112042 19848
rect 112668 19836 112674 19848
rect 112036 19808 112674 19836
rect 112036 19796 112042 19808
rect 112668 19796 112674 19808
rect 112726 19796 112732 19848
rect 114646 19796 114652 19848
rect 114704 19836 114710 19848
rect 115428 19836 115434 19848
rect 114704 19808 115434 19836
rect 114704 19796 114710 19808
rect 115428 19796 115434 19808
rect 115486 19796 115492 19848
rect 122806 19836 122834 19876
rect 132466 19876 150900 19904
rect 127434 19836 127440 19848
rect 122806 19808 127440 19836
rect 127434 19796 127440 19808
rect 127492 19796 127498 19848
rect 127894 19796 127900 19848
rect 127952 19836 127958 19848
rect 132466 19836 132494 19876
rect 150894 19864 150900 19876
rect 150952 19864 150958 19916
rect 152458 19864 152464 19916
rect 152516 19904 152522 19916
rect 153378 19904 153384 19916
rect 152516 19876 153384 19904
rect 152516 19864 152522 19876
rect 153378 19864 153384 19876
rect 153436 19864 153442 19916
rect 156782 19864 156788 19916
rect 156840 19904 156846 19916
rect 178126 19904 178132 19916
rect 156840 19876 178132 19904
rect 156840 19864 156846 19876
rect 178126 19864 178132 19876
rect 178184 19864 178190 19916
rect 127952 19808 132494 19836
rect 127952 19796 127958 19808
rect 150618 19796 150624 19848
rect 150676 19836 150682 19848
rect 152550 19836 152556 19848
rect 150676 19808 152556 19836
rect 150676 19796 150682 19808
rect 152550 19796 152556 19808
rect 152608 19796 152614 19848
rect 153746 19796 153752 19848
rect 153804 19836 153810 19848
rect 156506 19836 156512 19848
rect 153804 19808 156512 19836
rect 153804 19796 153810 19808
rect 156506 19796 156512 19808
rect 156564 19796 156570 19848
rect 156598 19796 156604 19848
rect 156656 19836 156662 19848
rect 211062 19836 211068 19848
rect 156656 19808 211068 19836
rect 156656 19796 156662 19808
rect 211062 19796 211068 19808
rect 211120 19796 211126 19848
rect 151170 19728 151176 19780
rect 151228 19768 151234 19780
rect 153010 19768 153016 19780
rect 151228 19740 153016 19768
rect 151228 19728 151234 19740
rect 153010 19728 153016 19740
rect 153068 19728 153074 19780
rect 155310 19728 155316 19780
rect 155368 19768 155374 19780
rect 155368 19740 157656 19768
rect 155368 19728 155374 19740
rect 104434 19700 104440 19712
rect 103486 19672 104440 19700
rect 81492 19660 81498 19672
rect 104434 19660 104440 19672
rect 104492 19660 104498 19712
rect 111150 19660 111156 19712
rect 111208 19700 111214 19712
rect 117406 19700 117412 19712
rect 111208 19672 117412 19700
rect 111208 19660 111214 19672
rect 117406 19660 117412 19672
rect 117464 19660 117470 19712
rect 149054 19660 149060 19712
rect 149112 19700 149118 19712
rect 152458 19700 152464 19712
rect 149112 19672 152464 19700
rect 149112 19660 149118 19672
rect 152458 19660 152464 19672
rect 152516 19660 152522 19712
rect 152550 19660 152556 19712
rect 152608 19700 152614 19712
rect 157242 19700 157248 19712
rect 152608 19672 157248 19700
rect 152608 19660 152614 19672
rect 157242 19660 157248 19672
rect 157300 19660 157306 19712
rect 157628 19700 157656 19740
rect 157702 19728 157708 19780
rect 157760 19768 157766 19780
rect 237374 19768 237380 19780
rect 157760 19740 237380 19768
rect 157760 19728 157766 19740
rect 237374 19728 237380 19740
rect 237432 19728 237438 19780
rect 247034 19700 247040 19712
rect 157628 19672 247040 19700
rect 247034 19660 247040 19672
rect 247092 19660 247098 19712
rect 16298 19592 16304 19644
rect 16356 19632 16362 19644
rect 21358 19632 21364 19644
rect 16356 19604 21364 19632
rect 16356 19592 16362 19604
rect 21358 19592 21364 19604
rect 21416 19592 21422 19644
rect 82814 19592 82820 19644
rect 82872 19632 82878 19644
rect 121546 19632 121552 19644
rect 82872 19604 121552 19632
rect 82872 19592 82878 19604
rect 121546 19592 121552 19604
rect 121604 19592 121610 19644
rect 122006 19592 122012 19644
rect 122064 19632 122070 19644
rect 126790 19632 126796 19644
rect 122064 19604 126796 19632
rect 122064 19592 122070 19604
rect 126790 19592 126796 19604
rect 126848 19592 126854 19644
rect 128446 19592 128452 19644
rect 128504 19632 128510 19644
rect 142614 19632 142620 19644
rect 128504 19604 142620 19632
rect 128504 19592 128510 19604
rect 142614 19592 142620 19604
rect 142672 19592 142678 19644
rect 150434 19592 150440 19644
rect 150492 19632 150498 19644
rect 154206 19632 154212 19644
rect 150492 19604 154212 19632
rect 150492 19592 150498 19604
rect 154206 19592 154212 19604
rect 154264 19592 154270 19644
rect 155954 19592 155960 19644
rect 156012 19632 156018 19644
rect 270402 19632 270408 19644
rect 156012 19604 270408 19632
rect 156012 19592 156018 19604
rect 270402 19592 270408 19604
rect 270460 19592 270466 19644
rect 102594 19524 102600 19576
rect 102652 19564 102658 19576
rect 131114 19564 131120 19576
rect 102652 19536 131120 19564
rect 102652 19524 102658 19536
rect 131114 19524 131120 19536
rect 131172 19524 131178 19576
rect 152182 19524 152188 19576
rect 152240 19564 152246 19576
rect 266354 19564 266360 19576
rect 152240 19536 266360 19564
rect 152240 19524 152246 19536
rect 266354 19524 266360 19536
rect 266412 19524 266418 19576
rect 103698 19456 103704 19508
rect 103756 19496 103762 19508
rect 148318 19496 148324 19508
rect 103756 19468 148324 19496
rect 103756 19456 103762 19468
rect 148318 19456 148324 19468
rect 148376 19456 148382 19508
rect 154574 19456 154580 19508
rect 154632 19496 154638 19508
rect 157702 19496 157708 19508
rect 154632 19468 157708 19496
rect 154632 19456 154638 19468
rect 157702 19456 157708 19468
rect 157760 19456 157766 19508
rect 157794 19456 157800 19508
rect 157852 19496 157858 19508
rect 460290 19496 460296 19508
rect 157852 19468 460296 19496
rect 157852 19456 157858 19468
rect 460290 19456 460296 19468
rect 460348 19456 460354 19508
rect 87966 19388 87972 19440
rect 88024 19428 88030 19440
rect 99190 19428 99196 19440
rect 88024 19400 99196 19428
rect 88024 19388 88030 19400
rect 99190 19388 99196 19400
rect 99248 19388 99254 19440
rect 112530 19388 112536 19440
rect 112588 19428 112594 19440
rect 437474 19428 437480 19440
rect 112588 19400 437480 19428
rect 112588 19388 112594 19400
rect 437474 19388 437480 19400
rect 437532 19388 437538 19440
rect 63402 19320 63408 19372
rect 63460 19360 63466 19372
rect 94222 19360 94228 19372
rect 63460 19332 94228 19360
rect 63460 19320 63466 19332
rect 94222 19320 94228 19332
rect 94280 19320 94286 19372
rect 96522 19320 96528 19372
rect 96580 19360 96586 19372
rect 102962 19360 102968 19372
rect 96580 19332 102968 19360
rect 96580 19320 96586 19332
rect 102962 19320 102968 19332
rect 103020 19320 103026 19372
rect 104802 19320 104808 19372
rect 104860 19360 104866 19372
rect 104860 19332 114554 19360
rect 104860 19320 104866 19332
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 81434 19292 81440 19304
rect 17644 19264 81440 19292
rect 17644 19252 17650 19264
rect 81434 19252 81440 19264
rect 81492 19252 81498 19304
rect 114526 19292 114554 19332
rect 118418 19320 118424 19372
rect 118476 19360 118482 19372
rect 121914 19360 121920 19372
rect 118476 19332 121920 19360
rect 118476 19320 118482 19332
rect 121914 19320 121920 19332
rect 121972 19320 121978 19372
rect 122098 19320 122104 19372
rect 122156 19360 122162 19372
rect 124950 19360 124956 19372
rect 122156 19332 124956 19360
rect 122156 19320 122162 19332
rect 124950 19320 124956 19332
rect 125008 19320 125014 19372
rect 127434 19320 127440 19372
rect 127492 19360 127498 19372
rect 513374 19360 513380 19372
rect 127492 19332 513380 19360
rect 127492 19320 127498 19332
rect 513374 19320 513380 19332
rect 513432 19320 513438 19372
rect 114526 19264 118694 19292
rect 18598 19184 18604 19236
rect 18656 19224 18662 19236
rect 23382 19224 23388 19236
rect 18656 19196 23388 19224
rect 18656 19184 18662 19196
rect 23382 19184 23388 19196
rect 23440 19184 23446 19236
rect 60090 19184 60096 19236
rect 60148 19224 60154 19236
rect 115290 19224 115296 19236
rect 60148 19196 115296 19224
rect 60148 19184 60154 19196
rect 115290 19184 115296 19196
rect 115348 19184 115354 19236
rect 118666 19224 118694 19264
rect 153654 19252 153660 19304
rect 153712 19292 153718 19304
rect 156046 19292 156052 19304
rect 153712 19264 156052 19292
rect 153712 19252 153718 19264
rect 156046 19252 156052 19264
rect 156104 19252 156110 19304
rect 222930 19252 222936 19304
rect 222988 19292 222994 19304
rect 226426 19292 226432 19304
rect 222988 19264 226432 19292
rect 222988 19252 222994 19264
rect 226426 19252 226432 19264
rect 226484 19252 226490 19304
rect 377398 19252 377404 19304
rect 377456 19292 377462 19304
rect 381906 19292 381912 19304
rect 377456 19264 381912 19292
rect 377456 19252 377462 19264
rect 381906 19252 381912 19264
rect 381964 19252 381970 19304
rect 150434 19224 150440 19236
rect 118666 19196 150440 19224
rect 150434 19184 150440 19196
rect 150492 19184 150498 19236
rect 154298 19184 154304 19236
rect 154356 19224 154362 19236
rect 154574 19224 154580 19236
rect 154356 19196 154580 19224
rect 154356 19184 154362 19196
rect 154574 19184 154580 19196
rect 154632 19184 154638 19236
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 69382 19156 69388 19168
rect 12124 19128 69388 19156
rect 12124 19116 12130 19128
rect 69382 19116 69388 19128
rect 69440 19116 69446 19168
rect 74994 19116 75000 19168
rect 75052 19156 75058 19168
rect 119338 19156 119344 19168
rect 75052 19128 119344 19156
rect 75052 19116 75058 19128
rect 119338 19116 119344 19128
rect 119396 19116 119402 19168
rect 121914 19116 121920 19168
rect 121972 19156 121978 19168
rect 124582 19156 124588 19168
rect 121972 19128 124588 19156
rect 121972 19116 121978 19128
rect 124582 19116 124588 19128
rect 124640 19116 124646 19168
rect 128170 19116 128176 19168
rect 128228 19156 128234 19168
rect 149054 19156 149060 19168
rect 128228 19128 149060 19156
rect 128228 19116 128234 19128
rect 149054 19116 149060 19128
rect 149112 19116 149118 19168
rect 62298 19048 62304 19100
rect 62356 19088 62362 19100
rect 62356 19060 103514 19088
rect 62356 19048 62362 19060
rect 18782 18980 18788 19032
rect 18840 19020 18846 19032
rect 84378 19020 84384 19032
rect 18840 18992 84384 19020
rect 18840 18980 18846 18992
rect 84378 18980 84384 18992
rect 84436 18980 84442 19032
rect 103486 19020 103514 19060
rect 121546 19048 121552 19100
rect 121604 19088 121610 19100
rect 129550 19088 129556 19100
rect 121604 19060 129556 19088
rect 121604 19048 121610 19060
rect 129550 19048 129556 19060
rect 129608 19048 129614 19100
rect 131114 19048 131120 19100
rect 131172 19088 131178 19100
rect 151078 19088 151084 19100
rect 131172 19060 151084 19088
rect 131172 19048 131178 19060
rect 151078 19048 151084 19060
rect 151136 19048 151142 19100
rect 247034 19048 247040 19100
rect 247092 19088 247098 19100
rect 260834 19088 260840 19100
rect 247092 19060 260840 19088
rect 247092 19048 247098 19060
rect 260834 19048 260840 19060
rect 260892 19048 260898 19100
rect 266354 19048 266360 19100
rect 266412 19088 266418 19100
rect 276014 19088 276020 19100
rect 266412 19060 276020 19088
rect 266412 19048 266418 19060
rect 276014 19048 276020 19060
rect 276072 19048 276078 19100
rect 122466 19020 122472 19032
rect 103486 18992 122472 19020
rect 122466 18980 122472 18992
rect 122524 18980 122530 19032
rect 124858 18980 124864 19032
rect 124916 19020 124922 19032
rect 128354 19020 128360 19032
rect 124916 18992 128360 19020
rect 124916 18980 124922 18992
rect 128354 18980 128360 18992
rect 128412 18980 128418 19032
rect 128538 18980 128544 19032
rect 128596 19020 128602 19032
rect 147674 19020 147680 19032
rect 128596 18992 147680 19020
rect 128596 18980 128602 18992
rect 147674 18980 147680 18992
rect 147732 18980 147738 19032
rect 149238 18980 149244 19032
rect 149296 19020 149302 19032
rect 151262 19020 151268 19032
rect 149296 18992 151268 19020
rect 149296 18980 149302 18992
rect 151262 18980 151268 18992
rect 151320 18980 151326 19032
rect 254026 18980 254032 19032
rect 254084 19020 254090 19032
rect 280430 19020 280436 19032
rect 254084 18992 280436 19020
rect 254084 18980 254090 18992
rect 280430 18980 280436 18992
rect 280488 18980 280494 19032
rect 19794 18912 19800 18964
rect 19852 18952 19858 18964
rect 86770 18952 86776 18964
rect 19852 18924 86776 18952
rect 19852 18912 19858 18924
rect 86770 18912 86776 18924
rect 86828 18912 86834 18964
rect 87690 18912 87696 18964
rect 87748 18952 87754 18964
rect 101122 18952 101128 18964
rect 87748 18924 101128 18952
rect 87748 18912 87754 18924
rect 101122 18912 101128 18924
rect 101180 18912 101186 18964
rect 111610 18912 111616 18964
rect 111668 18952 111674 18964
rect 152826 18952 152832 18964
rect 111668 18924 152832 18952
rect 111668 18912 111674 18924
rect 152826 18912 152832 18924
rect 152884 18912 152890 18964
rect 237374 18912 237380 18964
rect 237432 18952 237438 18964
rect 267826 18952 267832 18964
rect 237432 18924 267832 18952
rect 237432 18912 237438 18924
rect 267826 18912 267832 18924
rect 267884 18912 267890 18964
rect 6546 18844 6552 18896
rect 6604 18884 6610 18896
rect 15654 18884 15660 18896
rect 6604 18856 15660 18884
rect 6604 18844 6610 18856
rect 15654 18844 15660 18856
rect 15712 18844 15718 18896
rect 16206 18844 16212 18896
rect 16264 18884 16270 18896
rect 19058 18884 19064 18896
rect 16264 18856 19064 18884
rect 16264 18844 16270 18856
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 61194 18844 61200 18896
rect 61252 18884 61258 18896
rect 135346 18884 135352 18896
rect 61252 18856 135352 18884
rect 61252 18844 61258 18856
rect 135346 18844 135352 18856
rect 135404 18844 135410 18896
rect 151262 18844 151268 18896
rect 151320 18884 151326 18896
rect 155770 18884 155776 18896
rect 151320 18856 155776 18884
rect 151320 18844 151326 18856
rect 155770 18844 155776 18856
rect 155828 18844 155834 18896
rect 178126 18844 178132 18896
rect 178184 18884 178190 18896
rect 283374 18884 283380 18896
rect 178184 18856 283380 18884
rect 178184 18844 178190 18856
rect 283374 18844 283380 18856
rect 283432 18844 283438 18896
rect 336090 18844 336096 18896
rect 336148 18884 336154 18896
rect 381538 18884 381544 18896
rect 336148 18856 381544 18884
rect 336148 18844 336154 18856
rect 381538 18844 381544 18856
rect 381596 18844 381602 18896
rect 388346 18844 388352 18896
rect 388404 18884 388410 18896
rect 439222 18884 439228 18896
rect 388404 18856 439228 18884
rect 388404 18844 388410 18856
rect 439222 18844 439228 18856
rect 439280 18844 439286 18896
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 67174 18816 67180 18828
rect 11848 18788 67180 18816
rect 11848 18776 11854 18788
rect 67174 18776 67180 18788
rect 67232 18776 67238 18828
rect 73522 18776 73528 18828
rect 73580 18816 73586 18828
rect 215294 18816 215300 18828
rect 73580 18788 215300 18816
rect 73580 18776 73586 18788
rect 215294 18776 215300 18788
rect 215352 18776 215358 18828
rect 260742 18776 260748 18828
rect 260800 18816 260806 18828
rect 388438 18816 388444 18828
rect 260800 18788 388444 18816
rect 260800 18776 260806 18788
rect 388438 18776 388444 18788
rect 388496 18776 388502 18828
rect 403894 18776 403900 18828
rect 403952 18816 403958 18828
rect 470594 18816 470600 18828
rect 403952 18788 470600 18816
rect 403952 18776 403958 18788
rect 470594 18776 470600 18788
rect 470652 18776 470658 18828
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 15378 18748 15384 18760
rect 5132 18720 15384 18748
rect 5132 18708 5138 18720
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 64966 18748 64972 18760
rect 17552 18720 64972 18748
rect 17552 18708 17558 18720
rect 64966 18708 64972 18720
rect 65024 18708 65030 18760
rect 80514 18708 80520 18760
rect 80572 18748 80578 18760
rect 248506 18748 248512 18760
rect 80572 18720 248512 18748
rect 80572 18708 80578 18720
rect 248506 18708 248512 18720
rect 248564 18708 248570 18760
rect 270402 18708 270408 18760
rect 270460 18748 270466 18760
rect 408494 18748 408500 18760
rect 270460 18720 408500 18748
rect 270460 18708 270466 18720
rect 408494 18708 408500 18720
rect 408552 18708 408558 18760
rect 408586 18708 408592 18760
rect 408644 18748 408650 18760
rect 417418 18748 417424 18760
rect 408644 18720 417424 18748
rect 408644 18708 408650 18720
rect 417418 18708 417424 18720
rect 417476 18708 417482 18760
rect 4982 18640 4988 18692
rect 5040 18680 5046 18692
rect 15194 18680 15200 18692
rect 5040 18652 15200 18680
rect 5040 18640 5046 18652
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 16114 18640 16120 18692
rect 16172 18680 16178 18692
rect 35986 18680 35992 18692
rect 16172 18652 35992 18680
rect 16172 18640 16178 18652
rect 35986 18640 35992 18652
rect 36044 18640 36050 18692
rect 36170 18640 36176 18692
rect 36228 18680 36234 18692
rect 73798 18680 73804 18692
rect 36228 18652 73804 18680
rect 36228 18640 36234 18652
rect 73798 18640 73804 18652
rect 73856 18640 73862 18692
rect 82170 18640 82176 18692
rect 82228 18680 82234 18692
rect 270494 18680 270500 18692
rect 82228 18652 270500 18680
rect 82228 18640 82234 18652
rect 270494 18640 270500 18652
rect 270552 18640 270558 18692
rect 299382 18640 299388 18692
rect 299440 18680 299446 18692
rect 560294 18680 560300 18692
rect 299440 18652 560300 18680
rect 299440 18640 299446 18652
rect 560294 18640 560300 18652
rect 560352 18640 560358 18692
rect 2406 18572 2412 18624
rect 2464 18612 2470 18624
rect 2464 18584 2774 18612
rect 2464 18572 2470 18584
rect 2746 18476 2774 18584
rect 13354 18572 13360 18624
rect 13412 18612 13418 18624
rect 17678 18612 17684 18624
rect 13412 18584 17684 18612
rect 13412 18572 13418 18584
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 18690 18572 18696 18624
rect 18748 18612 18754 18624
rect 76098 18612 76104 18624
rect 18748 18584 31248 18612
rect 18748 18572 18754 18584
rect 17310 18504 17316 18556
rect 17368 18544 17374 18556
rect 31220 18544 31248 18584
rect 31726 18584 76104 18612
rect 31726 18544 31754 18584
rect 76098 18572 76104 18584
rect 76156 18572 76162 18624
rect 77754 18572 77760 18624
rect 77812 18612 77818 18624
rect 210050 18612 210056 18624
rect 77812 18584 210056 18612
rect 77812 18572 77818 18584
rect 210050 18572 210056 18584
rect 210108 18572 210114 18624
rect 211062 18572 211068 18624
rect 211120 18612 211126 18624
rect 502978 18612 502984 18624
rect 211120 18584 502984 18612
rect 211120 18572 211126 18584
rect 502978 18572 502984 18584
rect 503036 18572 503042 18624
rect 17368 18516 29684 18544
rect 31220 18516 31754 18544
rect 17368 18504 17374 18516
rect 18046 18476 18052 18488
rect 2746 18448 18052 18476
rect 18046 18436 18052 18448
rect 18104 18436 18110 18488
rect 19150 18436 19156 18488
rect 19208 18476 19214 18488
rect 29656 18476 29684 18516
rect 35802 18504 35808 18556
rect 35860 18544 35866 18556
rect 69934 18544 69940 18556
rect 35860 18516 69940 18544
rect 35860 18504 35866 18516
rect 69934 18504 69940 18516
rect 69992 18504 69998 18556
rect 129090 18504 129096 18556
rect 129148 18544 129154 18556
rect 146938 18544 146944 18556
rect 129148 18516 146944 18544
rect 129148 18504 129154 18516
rect 146938 18504 146944 18516
rect 146996 18504 147002 18556
rect 149146 18504 149152 18556
rect 149204 18544 149210 18556
rect 151906 18544 151912 18556
rect 149204 18516 151912 18544
rect 149204 18504 149210 18516
rect 151906 18504 151912 18516
rect 151964 18504 151970 18556
rect 33502 18476 33508 18488
rect 19208 18448 26234 18476
rect 29656 18448 33508 18476
rect 19208 18436 19214 18448
rect 26206 18408 26234 18448
rect 33502 18436 33508 18448
rect 33560 18436 33566 18488
rect 66438 18436 66444 18488
rect 66496 18476 66502 18488
rect 85390 18476 85396 18488
rect 66496 18448 85396 18476
rect 66496 18436 66502 18448
rect 85390 18436 85396 18448
rect 85448 18436 85454 18488
rect 100846 18436 100852 18488
rect 100904 18476 100910 18488
rect 101306 18476 101312 18488
rect 100904 18448 101312 18476
rect 100904 18436 100910 18448
rect 101306 18436 101312 18448
rect 101364 18436 101370 18488
rect 104986 18436 104992 18488
rect 105044 18476 105050 18488
rect 105170 18476 105176 18488
rect 105044 18448 105176 18476
rect 105044 18436 105050 18448
rect 105170 18436 105176 18448
rect 105228 18436 105234 18488
rect 150526 18436 150532 18488
rect 150584 18476 150590 18488
rect 154482 18476 154488 18488
rect 150584 18448 154488 18476
rect 150584 18436 150590 18448
rect 154482 18436 154488 18448
rect 154540 18436 154546 18488
rect 31662 18408 31668 18420
rect 26206 18380 31668 18408
rect 31662 18368 31668 18380
rect 31720 18368 31726 18420
rect 41598 18368 41604 18420
rect 41656 18408 41662 18420
rect 41782 18408 41788 18420
rect 41656 18380 41788 18408
rect 41656 18368 41662 18380
rect 41782 18368 41788 18380
rect 41840 18368 41846 18420
rect 42886 18368 42892 18420
rect 42944 18408 42950 18420
rect 43070 18408 43076 18420
rect 42944 18380 43076 18408
rect 42944 18368 42950 18380
rect 43070 18368 43076 18380
rect 43128 18368 43134 18420
rect 84930 18368 84936 18420
rect 84988 18408 84994 18420
rect 157426 18408 157432 18420
rect 84988 18380 157432 18408
rect 84988 18368 84994 18380
rect 157426 18368 157432 18380
rect 157484 18368 157490 18420
rect 10502 18300 10508 18352
rect 10560 18340 10566 18352
rect 68830 18340 68836 18352
rect 10560 18312 68836 18340
rect 10560 18300 10566 18312
rect 68830 18300 68836 18312
rect 68888 18300 68894 18352
rect 70578 18300 70584 18352
rect 70636 18340 70642 18352
rect 71222 18340 71228 18352
rect 70636 18312 71228 18340
rect 70636 18300 70642 18312
rect 71222 18300 71228 18312
rect 71280 18300 71286 18352
rect 79962 18300 79968 18352
rect 80020 18340 80026 18352
rect 116670 18340 116676 18352
rect 80020 18312 116676 18340
rect 80020 18300 80026 18312
rect 116670 18300 116676 18312
rect 116728 18300 116734 18352
rect 120074 18300 120080 18352
rect 120132 18340 120138 18352
rect 120718 18340 120724 18352
rect 120132 18312 120724 18340
rect 120132 18300 120138 18312
rect 120718 18300 120724 18312
rect 120776 18300 120782 18352
rect 123110 18300 123116 18352
rect 123168 18340 123174 18352
rect 128446 18340 128452 18352
rect 123168 18312 128452 18340
rect 123168 18300 123174 18312
rect 128446 18300 128452 18312
rect 128504 18300 128510 18352
rect 149054 18300 149060 18352
rect 149112 18340 149118 18352
rect 321554 18340 321560 18352
rect 149112 18312 321560 18340
rect 149112 18300 149118 18312
rect 321554 18300 321560 18312
rect 321612 18300 321618 18352
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 65518 18272 65524 18284
rect 16448 18244 65524 18272
rect 16448 18232 16454 18244
rect 65518 18232 65524 18244
rect 65576 18232 65582 18284
rect 98086 18232 98092 18284
rect 98144 18272 98150 18284
rect 99006 18272 99012 18284
rect 98144 18244 99012 18272
rect 98144 18232 98150 18244
rect 99006 18232 99012 18244
rect 99064 18232 99070 18284
rect 100846 18232 100852 18284
rect 100904 18272 100910 18284
rect 101398 18272 101404 18284
rect 100904 18244 101404 18272
rect 100904 18232 100910 18244
rect 101398 18232 101404 18244
rect 101456 18232 101462 18284
rect 102134 18232 102140 18284
rect 102192 18272 102198 18284
rect 113818 18272 113824 18284
rect 102192 18244 113824 18272
rect 102192 18232 102198 18244
rect 113818 18232 113824 18244
rect 113876 18232 113882 18284
rect 120994 18232 121000 18284
rect 121052 18272 121058 18284
rect 128354 18272 128360 18284
rect 121052 18244 128360 18272
rect 121052 18232 121058 18244
rect 128354 18232 128360 18244
rect 128412 18232 128418 18284
rect 153010 18232 153016 18284
rect 153068 18272 153074 18284
rect 239582 18272 239588 18284
rect 153068 18244 239588 18272
rect 153068 18232 153074 18244
rect 239582 18232 239588 18244
rect 239640 18232 239646 18284
rect 7834 18164 7840 18216
rect 7892 18204 7898 18216
rect 63402 18204 63408 18216
rect 7892 18176 63408 18204
rect 7892 18164 7898 18176
rect 63402 18164 63408 18176
rect 63460 18164 63466 18216
rect 95142 18164 95148 18216
rect 95200 18204 95206 18216
rect 187602 18204 187608 18216
rect 95200 18176 187608 18204
rect 95200 18164 95206 18176
rect 187602 18164 187608 18176
rect 187660 18164 187666 18216
rect 14642 18096 14648 18148
rect 14700 18136 14706 18148
rect 17770 18136 17776 18148
rect 14700 18108 17776 18136
rect 14700 18096 14706 18108
rect 17770 18096 17776 18108
rect 17828 18096 17834 18148
rect 43162 18096 43168 18148
rect 43220 18136 43226 18148
rect 43622 18136 43628 18148
rect 43220 18108 43628 18136
rect 43220 18096 43226 18108
rect 43622 18096 43628 18108
rect 43680 18096 43686 18148
rect 85482 18096 85488 18148
rect 85540 18136 85546 18148
rect 112438 18136 112444 18148
rect 85540 18108 112444 18136
rect 85540 18096 85546 18108
rect 112438 18096 112444 18108
rect 112496 18096 112502 18148
rect 116026 18096 116032 18148
rect 116084 18136 116090 18148
rect 124306 18136 124312 18148
rect 116084 18108 124312 18136
rect 116084 18096 116090 18108
rect 124306 18096 124312 18108
rect 124364 18096 124370 18148
rect 147766 18096 147772 18148
rect 147824 18136 147830 18148
rect 150618 18136 150624 18148
rect 147824 18108 150624 18136
rect 147824 18096 147830 18108
rect 150618 18096 150624 18108
rect 150676 18096 150682 18148
rect 150894 18096 150900 18148
rect 150952 18136 150958 18148
rect 152182 18136 152188 18148
rect 150952 18108 152188 18136
rect 150952 18096 150958 18108
rect 152182 18096 152188 18108
rect 152240 18096 152246 18148
rect 154206 18096 154212 18148
rect 154264 18136 154270 18148
rect 155862 18136 155868 18148
rect 154264 18108 155868 18136
rect 154264 18096 154270 18108
rect 155862 18096 155868 18108
rect 155920 18096 155926 18148
rect 158438 18096 158444 18148
rect 158496 18136 158502 18148
rect 263134 18136 263140 18148
rect 158496 18108 263140 18136
rect 158496 18096 158502 18108
rect 263134 18096 263140 18108
rect 263192 18096 263198 18148
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 16942 18068 16948 18080
rect 14608 18040 16948 18068
rect 14608 18028 14614 18040
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 43070 18028 43076 18080
rect 43128 18068 43134 18080
rect 43438 18068 43444 18080
rect 43128 18040 43444 18068
rect 43128 18028 43134 18040
rect 43438 18028 43444 18040
rect 43496 18028 43502 18080
rect 85758 18028 85764 18080
rect 85816 18068 85822 18080
rect 87966 18068 87972 18080
rect 85816 18040 87972 18068
rect 85816 18028 85822 18040
rect 87966 18028 87972 18040
rect 88024 18028 88030 18080
rect 244550 18068 244556 18080
rect 103486 18040 244556 18068
rect 14458 17960 14464 18012
rect 14516 18000 14522 18012
rect 16758 18000 16764 18012
rect 14516 17972 16764 18000
rect 14516 17960 14522 17972
rect 16758 17960 16764 17972
rect 16816 17960 16822 18012
rect 78646 17972 91140 18000
rect 10594 17892 10600 17944
rect 10652 17932 10658 17944
rect 13262 17932 13268 17944
rect 10652 17904 13268 17932
rect 10652 17892 10658 17904
rect 13262 17892 13268 17904
rect 13320 17892 13326 17944
rect 19978 17892 19984 17944
rect 20036 17932 20042 17944
rect 23106 17932 23112 17944
rect 20036 17904 23112 17932
rect 20036 17892 20042 17904
rect 23106 17892 23112 17904
rect 23164 17892 23170 17944
rect 40770 17892 40776 17944
rect 40828 17932 40834 17944
rect 42058 17932 42064 17944
rect 40828 17904 42064 17932
rect 40828 17892 40834 17904
rect 42058 17892 42064 17904
rect 42116 17892 42122 17944
rect 45554 17892 45560 17944
rect 45612 17932 45618 17944
rect 47118 17932 47124 17944
rect 45612 17904 47124 17932
rect 45612 17892 45618 17904
rect 47118 17892 47124 17904
rect 47176 17892 47182 17944
rect 48498 17892 48504 17944
rect 48556 17932 48562 17944
rect 50706 17932 50712 17944
rect 48556 17904 50712 17932
rect 48556 17892 48562 17904
rect 50706 17892 50712 17904
rect 50764 17892 50770 17944
rect 52178 17892 52184 17944
rect 52236 17932 52242 17944
rect 52454 17932 52460 17944
rect 52236 17904 52460 17932
rect 52236 17892 52242 17904
rect 52454 17892 52460 17904
rect 52512 17892 52518 17944
rect 60642 17892 60648 17944
rect 60700 17932 60706 17944
rect 63310 17932 63316 17944
rect 60700 17904 63316 17932
rect 60700 17892 60706 17904
rect 63310 17892 63316 17904
rect 63368 17892 63374 17944
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 13354 17864 13360 17876
rect 9456 17836 13360 17864
rect 9456 17824 9462 17836
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 67726 17864 67732 17876
rect 13504 17836 67732 17864
rect 13504 17824 13510 17836
rect 67726 17824 67732 17836
rect 67784 17824 67790 17876
rect 6638 17756 6644 17808
rect 6696 17796 6702 17808
rect 6696 17768 11008 17796
rect 6696 17756 6702 17768
rect 3510 17688 3516 17740
rect 3568 17728 3574 17740
rect 3568 17700 10916 17728
rect 3568 17688 3574 17700
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 10888 17592 10916 17700
rect 10980 17660 11008 17768
rect 12158 17756 12164 17808
rect 12216 17796 12222 17808
rect 66622 17796 66628 17808
rect 12216 17768 66628 17796
rect 12216 17756 12222 17768
rect 66622 17756 66628 17768
rect 66680 17756 66686 17808
rect 12250 17688 12256 17740
rect 12308 17728 12314 17740
rect 66070 17728 66076 17740
rect 12308 17700 66076 17728
rect 12308 17688 12314 17700
rect 66070 17688 66076 17700
rect 66128 17688 66134 17740
rect 67726 17688 67732 17740
rect 67784 17728 67790 17740
rect 78646 17728 78674 17972
rect 80330 17892 80336 17944
rect 80388 17932 80394 17944
rect 81434 17932 81440 17944
rect 80388 17904 81440 17932
rect 80388 17892 80394 17904
rect 81434 17892 81440 17904
rect 81492 17892 81498 17944
rect 86770 17892 86776 17944
rect 86828 17932 86834 17944
rect 90358 17932 90364 17944
rect 86828 17904 90364 17932
rect 86828 17892 86834 17904
rect 90358 17892 90364 17904
rect 90416 17892 90422 17944
rect 91112 17932 91140 17972
rect 94590 17932 94596 17944
rect 91112 17904 94596 17932
rect 94590 17892 94596 17904
rect 94648 17892 94654 17944
rect 96706 17892 96712 17944
rect 96764 17932 96770 17944
rect 97902 17932 97908 17944
rect 96764 17904 97908 17932
rect 96764 17892 96770 17904
rect 97902 17892 97908 17904
rect 97960 17892 97966 17944
rect 98730 17892 98736 17944
rect 98788 17932 98794 17944
rect 100110 17932 100116 17944
rect 98788 17904 100116 17932
rect 98788 17892 98794 17904
rect 100110 17892 100116 17904
rect 100168 17892 100174 17944
rect 82722 17824 82728 17876
rect 82780 17864 82786 17876
rect 102134 17864 102140 17876
rect 82780 17836 102140 17864
rect 82780 17824 82786 17836
rect 102134 17824 102140 17836
rect 102192 17824 102198 17876
rect 89714 17756 89720 17808
rect 89772 17796 89778 17808
rect 91462 17796 91468 17808
rect 89772 17768 91468 17796
rect 89772 17756 89778 17768
rect 91462 17756 91468 17768
rect 91520 17756 91526 17808
rect 92566 17756 92572 17808
rect 92624 17796 92630 17808
rect 93118 17796 93124 17808
rect 92624 17768 93124 17796
rect 92624 17756 92630 17768
rect 93118 17756 93124 17768
rect 93176 17756 93182 17808
rect 103486 17796 103514 18040
rect 244550 18028 244556 18040
rect 244608 18028 244614 18080
rect 109006 17972 112024 18000
rect 108298 17892 108304 17944
rect 108356 17932 108362 17944
rect 109006 17932 109034 17972
rect 108356 17904 109034 17932
rect 108356 17892 108362 17904
rect 107378 17824 107384 17876
rect 107436 17864 107442 17876
rect 109586 17864 109592 17876
rect 107436 17836 109592 17864
rect 107436 17824 107442 17836
rect 109586 17824 109592 17836
rect 109644 17824 109650 17876
rect 110506 17824 110512 17876
rect 110564 17864 110570 17876
rect 111886 17864 111892 17876
rect 110564 17836 111892 17864
rect 110564 17824 110570 17836
rect 111886 17824 111892 17836
rect 111944 17824 111950 17876
rect 111996 17864 112024 17972
rect 113818 17960 113824 18012
rect 113876 18000 113882 18012
rect 120718 18000 120724 18012
rect 113876 17972 120724 18000
rect 113876 17960 113882 17972
rect 120718 17960 120724 17972
rect 120776 17960 120782 18012
rect 121546 17960 121552 18012
rect 121604 18000 121610 18012
rect 124030 18000 124036 18012
rect 121604 17972 124036 18000
rect 121604 17960 121610 17972
rect 124030 17960 124036 17972
rect 124088 17960 124094 18012
rect 136082 17960 136088 18012
rect 136140 18000 136146 18012
rect 146202 18000 146208 18012
rect 136140 17972 146208 18000
rect 136140 17960 136146 17972
rect 146202 17960 146208 17972
rect 146260 17960 146266 18012
rect 146956 17972 149100 18000
rect 118234 17892 118240 17944
rect 118292 17932 118298 17944
rect 121362 17932 121368 17944
rect 118292 17904 121368 17932
rect 118292 17892 118298 17904
rect 121362 17892 121368 17904
rect 121420 17892 121426 17944
rect 123202 17892 123208 17944
rect 123260 17932 123266 17944
rect 126514 17932 126520 17944
rect 123260 17904 126520 17932
rect 123260 17892 123266 17904
rect 126514 17892 126520 17904
rect 126572 17892 126578 17944
rect 137278 17892 137284 17944
rect 137336 17932 137342 17944
rect 146956 17932 146984 17972
rect 137336 17904 146984 17932
rect 149072 17932 149100 17972
rect 151170 17960 151176 18012
rect 151228 18000 151234 18012
rect 151446 18000 151452 18012
rect 151228 17972 151452 18000
rect 151228 17960 151234 17972
rect 151446 17960 151452 17972
rect 151504 17960 151510 18012
rect 160186 18000 160192 18012
rect 155972 17972 160192 18000
rect 151906 17932 151912 17944
rect 149072 17904 151912 17932
rect 137336 17892 137342 17904
rect 151906 17892 151912 17904
rect 151964 17892 151970 17944
rect 151998 17892 152004 17944
rect 152056 17932 152062 17944
rect 155972 17932 156000 17972
rect 160186 17960 160192 17972
rect 160244 17960 160250 18012
rect 152056 17904 156000 17932
rect 152056 17892 152062 17904
rect 424962 17892 424968 17944
rect 425020 17932 425026 17944
rect 431310 17932 431316 17944
rect 425020 17904 431316 17932
rect 425020 17892 425026 17904
rect 431310 17892 431316 17904
rect 431368 17892 431374 17944
rect 442258 17892 442264 17944
rect 442316 17932 442322 17944
rect 445478 17932 445484 17944
rect 442316 17904 445484 17932
rect 442316 17892 442322 17904
rect 445478 17892 445484 17904
rect 445536 17892 445542 17944
rect 471330 17892 471336 17944
rect 471388 17932 471394 17944
rect 473998 17932 474004 17944
rect 471388 17904 474004 17932
rect 471388 17892 471394 17904
rect 473998 17892 474004 17904
rect 474056 17892 474062 17944
rect 116578 17864 116584 17876
rect 111996 17836 116584 17864
rect 116578 17824 116584 17836
rect 116636 17824 116642 17876
rect 117866 17824 117872 17876
rect 117924 17864 117930 17876
rect 121270 17864 121276 17876
rect 117924 17836 121276 17864
rect 117924 17824 117930 17836
rect 121270 17824 121276 17836
rect 121328 17824 121334 17876
rect 143442 17824 143448 17876
rect 143500 17864 143506 17876
rect 149054 17864 149060 17876
rect 143500 17836 149060 17864
rect 143500 17824 143506 17836
rect 149054 17824 149060 17836
rect 149112 17824 149118 17876
rect 471422 17824 471428 17876
rect 471480 17864 471486 17876
rect 475378 17864 475384 17876
rect 471480 17836 475384 17864
rect 471480 17824 471486 17836
rect 475378 17824 475384 17836
rect 475436 17824 475442 17876
rect 93826 17768 103514 17796
rect 67784 17700 78674 17728
rect 67784 17688 67790 17700
rect 88058 17688 88064 17740
rect 88116 17728 88122 17740
rect 91554 17728 91560 17740
rect 88116 17700 91560 17728
rect 88116 17688 88122 17700
rect 91554 17688 91560 17700
rect 91612 17688 91618 17740
rect 18230 17660 18236 17672
rect 10980 17632 18236 17660
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 68278 17660 68284 17672
rect 23532 17632 68284 17660
rect 23532 17620 23538 17632
rect 68278 17620 68284 17632
rect 68336 17620 68342 17672
rect 68370 17620 68376 17672
rect 68428 17660 68434 17672
rect 68428 17632 76880 17660
rect 68428 17620 68434 17632
rect 36170 17592 36176 17604
rect 9272 17564 10824 17592
rect 10888 17564 36176 17592
rect 9272 17552 9278 17564
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 10686 17524 10692 17536
rect 7708 17496 10692 17524
rect 7708 17484 7714 17496
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 10796 17524 10824 17564
rect 36170 17552 36176 17564
rect 36228 17552 36234 17604
rect 40034 17552 40040 17604
rect 40092 17592 40098 17604
rect 42702 17592 42708 17604
rect 40092 17564 42708 17592
rect 40092 17552 40098 17564
rect 42702 17552 42708 17564
rect 42760 17552 42766 17604
rect 43346 17552 43352 17604
rect 43404 17592 43410 17604
rect 43404 17564 45554 17592
rect 43404 17552 43410 17564
rect 24854 17524 24860 17536
rect 10796 17496 24860 17524
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 27706 17484 27712 17536
rect 27764 17524 27770 17536
rect 44450 17524 44456 17536
rect 27764 17496 44456 17524
rect 27764 17484 27770 17496
rect 44450 17484 44456 17496
rect 44508 17484 44514 17536
rect 45526 17524 45554 17564
rect 51258 17552 51264 17604
rect 51316 17592 51322 17604
rect 53098 17592 53104 17604
rect 51316 17564 53104 17592
rect 51316 17552 51322 17564
rect 53098 17552 53104 17564
rect 53156 17552 53162 17604
rect 57514 17552 57520 17604
rect 57572 17592 57578 17604
rect 62022 17592 62028 17604
rect 57572 17564 62028 17592
rect 57572 17552 57578 17564
rect 62022 17552 62028 17564
rect 62080 17552 62086 17604
rect 63954 17552 63960 17604
rect 64012 17592 64018 17604
rect 66070 17592 66076 17604
rect 64012 17564 66076 17592
rect 64012 17552 64018 17564
rect 66070 17552 66076 17564
rect 66128 17552 66134 17604
rect 69290 17552 69296 17604
rect 69348 17592 69354 17604
rect 76852 17592 76880 17632
rect 77018 17620 77024 17672
rect 77076 17660 77082 17672
rect 79410 17660 79416 17672
rect 77076 17632 79416 17660
rect 77076 17620 77082 17632
rect 79410 17620 79416 17632
rect 79468 17620 79474 17672
rect 86586 17620 86592 17672
rect 86644 17660 86650 17672
rect 93118 17660 93124 17672
rect 86644 17632 93124 17660
rect 86644 17620 86650 17632
rect 93118 17620 93124 17632
rect 93176 17620 93182 17672
rect 79134 17592 79140 17604
rect 69348 17564 75408 17592
rect 76852 17564 79140 17592
rect 69348 17552 69354 17564
rect 62942 17524 62948 17536
rect 45526 17496 62948 17524
rect 62942 17484 62948 17496
rect 63000 17484 63006 17536
rect 65518 17484 65524 17536
rect 65576 17524 65582 17536
rect 75178 17524 75184 17536
rect 65576 17496 75184 17524
rect 65576 17484 65582 17496
rect 75178 17484 75184 17496
rect 75236 17484 75242 17536
rect 2222 17416 2228 17468
rect 2280 17456 2286 17468
rect 18138 17456 18144 17468
rect 2280 17428 18144 17456
rect 2280 17416 2286 17428
rect 18138 17416 18144 17428
rect 18196 17416 18202 17468
rect 19334 17416 19340 17468
rect 19392 17456 19398 17468
rect 42978 17456 42984 17468
rect 19392 17428 42984 17456
rect 19392 17416 19398 17428
rect 42978 17416 42984 17428
rect 43036 17416 43042 17468
rect 50338 17416 50344 17468
rect 50396 17456 50402 17468
rect 51810 17456 51816 17468
rect 50396 17428 51816 17456
rect 50396 17416 50402 17428
rect 51810 17416 51816 17428
rect 51868 17416 51874 17468
rect 52730 17416 52736 17468
rect 52788 17456 52794 17468
rect 73890 17456 73896 17468
rect 52788 17428 73896 17456
rect 52788 17416 52794 17428
rect 73890 17416 73896 17428
rect 73948 17416 73954 17468
rect 75380 17456 75408 17564
rect 79134 17552 79140 17564
rect 79192 17552 79198 17604
rect 87506 17552 87512 17604
rect 87564 17592 87570 17604
rect 90082 17592 90088 17604
rect 87564 17564 90088 17592
rect 87564 17552 87570 17564
rect 90082 17552 90088 17564
rect 90140 17552 90146 17604
rect 93826 17592 93854 17768
rect 104250 17756 104256 17808
rect 104308 17796 104314 17808
rect 108390 17796 108396 17808
rect 104308 17768 108396 17796
rect 104308 17756 104314 17768
rect 108390 17756 108396 17768
rect 108448 17756 108454 17808
rect 294598 17796 294604 17808
rect 109006 17768 294604 17796
rect 109006 17740 109034 17768
rect 294598 17756 294604 17768
rect 294656 17756 294662 17808
rect 322750 17796 322756 17808
rect 316006 17768 322756 17796
rect 97902 17688 97908 17740
rect 97960 17728 97966 17740
rect 107746 17728 107752 17740
rect 97960 17700 107752 17728
rect 97960 17688 97966 17700
rect 107746 17688 107752 17700
rect 107804 17688 107810 17740
rect 108942 17688 108948 17740
rect 109000 17700 109034 17740
rect 109000 17688 109006 17700
rect 109126 17688 109132 17740
rect 109184 17728 109190 17740
rect 113082 17728 113088 17740
rect 109184 17700 113088 17728
rect 109184 17688 109190 17700
rect 113082 17688 113088 17700
rect 113140 17688 113146 17740
rect 113726 17688 113732 17740
rect 113784 17728 113790 17740
rect 316006 17728 316034 17768
rect 322750 17756 322756 17768
rect 322808 17756 322814 17808
rect 113784 17700 316034 17728
rect 113784 17688 113790 17700
rect 321554 17688 321560 17740
rect 321612 17728 321618 17740
rect 373258 17728 373264 17740
rect 321612 17700 373264 17728
rect 321612 17688 321618 17700
rect 373258 17688 373264 17700
rect 373316 17688 373322 17740
rect 99466 17620 99472 17672
rect 99524 17660 99530 17672
rect 102318 17660 102324 17672
rect 99524 17632 102324 17660
rect 99524 17620 99530 17632
rect 102318 17620 102324 17632
rect 102376 17620 102382 17672
rect 212810 17660 212816 17672
rect 105464 17632 212816 17660
rect 92768 17564 93854 17592
rect 81986 17484 81992 17536
rect 82044 17524 82050 17536
rect 89254 17524 89260 17536
rect 82044 17496 89260 17524
rect 82044 17484 82050 17496
rect 89254 17484 89260 17496
rect 89312 17484 89318 17536
rect 82170 17456 82176 17468
rect 75380 17428 82176 17456
rect 82170 17416 82176 17428
rect 82228 17416 82234 17468
rect 84286 17416 84292 17468
rect 84344 17456 84350 17468
rect 92768 17456 92796 17564
rect 94130 17552 94136 17604
rect 94188 17592 94194 17604
rect 97074 17592 97080 17604
rect 94188 17564 97080 17592
rect 94188 17552 94194 17564
rect 97074 17552 97080 17564
rect 97132 17552 97138 17604
rect 97258 17552 97264 17604
rect 97316 17592 97322 17604
rect 97316 17564 99420 17592
rect 97316 17552 97322 17564
rect 92842 17484 92848 17536
rect 92900 17524 92906 17536
rect 99282 17524 99288 17536
rect 92900 17496 99288 17524
rect 92900 17484 92906 17496
rect 99282 17484 99288 17496
rect 99340 17484 99346 17536
rect 99392 17524 99420 17564
rect 101122 17552 101128 17604
rect 101180 17592 101186 17604
rect 105354 17592 105360 17604
rect 101180 17564 105360 17592
rect 101180 17552 101186 17564
rect 105354 17552 105360 17564
rect 105412 17552 105418 17604
rect 103054 17524 103060 17536
rect 99392 17496 103060 17524
rect 103054 17484 103060 17496
rect 103112 17484 103118 17536
rect 103422 17484 103428 17536
rect 103480 17524 103486 17536
rect 105464 17524 105492 17632
rect 212810 17620 212816 17632
rect 212868 17620 212874 17672
rect 239582 17620 239588 17672
rect 239640 17660 239646 17672
rect 477402 17660 477408 17672
rect 239640 17632 477408 17660
rect 239640 17620 239646 17632
rect 477402 17620 477408 17632
rect 477460 17620 477466 17672
rect 105722 17552 105728 17604
rect 105780 17592 105786 17604
rect 113358 17592 113364 17604
rect 105780 17564 113364 17592
rect 105780 17552 105786 17564
rect 113358 17552 113364 17564
rect 113416 17552 113422 17604
rect 114002 17552 114008 17604
rect 114060 17592 114066 17604
rect 372614 17592 372620 17604
rect 114060 17564 372620 17592
rect 114060 17552 114066 17564
rect 372614 17552 372620 17564
rect 372672 17552 372678 17604
rect 407022 17552 407028 17604
rect 407080 17592 407086 17604
rect 420914 17592 420920 17604
rect 407080 17564 420920 17592
rect 407080 17552 407086 17564
rect 420914 17552 420920 17564
rect 420972 17552 420978 17604
rect 421006 17552 421012 17604
rect 421064 17592 421070 17604
rect 427630 17592 427636 17604
rect 421064 17564 427636 17592
rect 421064 17552 421070 17564
rect 427630 17552 427636 17564
rect 427688 17552 427694 17604
rect 431218 17552 431224 17604
rect 431276 17592 431282 17604
rect 436002 17592 436008 17604
rect 431276 17564 436008 17592
rect 431276 17552 431282 17564
rect 436002 17552 436008 17564
rect 436060 17552 436066 17604
rect 103480 17496 105492 17524
rect 103480 17484 103486 17496
rect 106826 17484 106832 17536
rect 106884 17524 106890 17536
rect 378042 17524 378048 17536
rect 106884 17496 113864 17524
rect 106884 17484 106890 17496
rect 84344 17428 92796 17456
rect 84344 17416 84350 17428
rect 94130 17416 94136 17468
rect 94188 17456 94194 17468
rect 97534 17456 97540 17468
rect 94188 17428 97540 17456
rect 94188 17416 94194 17428
rect 97534 17416 97540 17428
rect 97592 17416 97598 17468
rect 103606 17416 103612 17468
rect 103664 17456 103670 17468
rect 109678 17456 109684 17468
rect 103664 17428 109684 17456
rect 103664 17416 103670 17428
rect 109678 17416 109684 17428
rect 109736 17416 109742 17468
rect 110138 17416 110144 17468
rect 110196 17456 110202 17468
rect 113726 17456 113732 17468
rect 110196 17428 113732 17456
rect 110196 17416 110202 17428
rect 113726 17416 113732 17428
rect 113784 17416 113790 17468
rect 113836 17456 113864 17496
rect 114112 17496 378048 17524
rect 114112 17456 114140 17496
rect 378042 17484 378048 17496
rect 378100 17484 378106 17536
rect 381630 17484 381636 17536
rect 381688 17524 381694 17536
rect 439406 17524 439412 17536
rect 381688 17496 439412 17524
rect 381688 17484 381694 17496
rect 439406 17484 439412 17496
rect 439464 17484 439470 17536
rect 113836 17428 114140 17456
rect 117682 17416 117688 17468
rect 117740 17456 117746 17468
rect 119522 17456 119528 17468
rect 117740 17428 119528 17456
rect 117740 17416 117746 17428
rect 119522 17416 119528 17428
rect 119580 17416 119586 17468
rect 120442 17416 120448 17468
rect 120500 17456 120506 17468
rect 122282 17456 122288 17468
rect 120500 17428 122288 17456
rect 120500 17416 120506 17428
rect 122282 17416 122288 17428
rect 122340 17416 122346 17468
rect 122374 17416 122380 17468
rect 122432 17456 122438 17468
rect 412634 17456 412640 17468
rect 122432 17428 412640 17456
rect 122432 17416 122438 17428
rect 412634 17416 412640 17428
rect 412692 17416 412698 17468
rect 435358 17416 435364 17468
rect 435416 17456 435422 17468
rect 448698 17456 448704 17468
rect 435416 17428 448704 17456
rect 435416 17416 435422 17428
rect 448698 17416 448704 17428
rect 448756 17416 448762 17468
rect 842 17348 848 17400
rect 900 17388 906 17400
rect 13446 17388 13452 17400
rect 900 17360 13452 17388
rect 900 17348 906 17360
rect 13446 17348 13452 17360
rect 13504 17348 13510 17400
rect 15562 17348 15568 17400
rect 15620 17388 15626 17400
rect 42334 17388 42340 17400
rect 15620 17360 42340 17388
rect 15620 17348 15626 17360
rect 42334 17348 42340 17360
rect 42392 17348 42398 17400
rect 45738 17348 45744 17400
rect 45796 17388 45802 17400
rect 65886 17388 65892 17400
rect 45796 17360 65892 17388
rect 45796 17348 45802 17360
rect 65886 17348 65892 17360
rect 65944 17348 65950 17400
rect 66254 17348 66260 17400
rect 66312 17388 66318 17400
rect 71590 17388 71596 17400
rect 66312 17360 71596 17388
rect 66312 17348 66318 17360
rect 71590 17348 71596 17360
rect 71648 17348 71654 17400
rect 75086 17348 75092 17400
rect 75144 17388 75150 17400
rect 80698 17388 80704 17400
rect 75144 17360 80704 17388
rect 75144 17348 75150 17360
rect 80698 17348 80704 17360
rect 80756 17348 80762 17400
rect 81066 17348 81072 17400
rect 81124 17388 81130 17400
rect 87598 17388 87604 17400
rect 81124 17360 87604 17388
rect 81124 17348 81130 17360
rect 87598 17348 87604 17360
rect 87656 17348 87662 17400
rect 90726 17348 90732 17400
rect 90784 17388 90790 17400
rect 97258 17388 97264 17400
rect 90784 17360 97264 17388
rect 90784 17348 90790 17360
rect 97258 17348 97264 17360
rect 97316 17348 97322 17400
rect 97350 17348 97356 17400
rect 97408 17388 97414 17400
rect 111334 17388 111340 17400
rect 97408 17360 111340 17388
rect 97408 17348 97414 17360
rect 111334 17348 111340 17360
rect 111392 17348 111398 17400
rect 113358 17348 113364 17400
rect 113416 17388 113422 17400
rect 422386 17388 422392 17400
rect 113416 17360 422392 17388
rect 113416 17348 113422 17360
rect 422386 17348 422392 17360
rect 422444 17348 422450 17400
rect 426802 17348 426808 17400
rect 426860 17388 426866 17400
rect 454770 17388 454776 17400
rect 426860 17360 454776 17388
rect 426860 17348 426866 17360
rect 454770 17348 454776 17360
rect 454828 17348 454834 17400
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 41414 17320 41420 17332
rect 9732 17292 41420 17320
rect 9732 17280 9738 17292
rect 41414 17280 41420 17292
rect 41472 17280 41478 17332
rect 43438 17280 43444 17332
rect 43496 17320 43502 17332
rect 44910 17320 44916 17332
rect 43496 17292 44916 17320
rect 43496 17280 43502 17292
rect 44910 17280 44916 17292
rect 44968 17280 44974 17332
rect 47946 17280 47952 17332
rect 48004 17320 48010 17332
rect 50338 17320 50344 17332
rect 48004 17292 50344 17320
rect 48004 17280 48010 17292
rect 50338 17280 50344 17292
rect 50396 17280 50402 17332
rect 54938 17280 54944 17332
rect 54996 17320 55002 17332
rect 61378 17320 61384 17332
rect 54996 17292 61384 17320
rect 54996 17280 55002 17292
rect 61378 17280 61384 17292
rect 61436 17280 61442 17332
rect 61838 17280 61844 17332
rect 61896 17320 61902 17332
rect 99190 17320 99196 17332
rect 61896 17292 99196 17320
rect 61896 17280 61902 17292
rect 99190 17280 99196 17292
rect 99248 17280 99254 17332
rect 100018 17280 100024 17332
rect 100076 17320 100082 17332
rect 109770 17320 109776 17332
rect 100076 17292 109776 17320
rect 100076 17280 100082 17292
rect 109770 17280 109776 17292
rect 109828 17280 109834 17332
rect 112346 17280 112352 17332
rect 112404 17320 112410 17332
rect 438118 17320 438124 17332
rect 112404 17292 438124 17320
rect 112404 17280 112410 17292
rect 438118 17280 438124 17292
rect 438176 17280 438182 17332
rect 36538 17212 36544 17264
rect 36596 17252 36602 17264
rect 45094 17252 45100 17264
rect 36596 17224 45100 17252
rect 36596 17212 36602 17224
rect 45094 17212 45100 17224
rect 45152 17212 45158 17264
rect 48222 17212 48228 17264
rect 48280 17252 48286 17264
rect 52730 17252 52736 17264
rect 48280 17224 52736 17252
rect 48280 17212 48286 17224
rect 52730 17212 52736 17224
rect 52788 17212 52794 17264
rect 59998 17252 60004 17264
rect 55186 17224 60004 17252
rect 2314 17144 2320 17196
rect 2372 17184 2378 17196
rect 8938 17184 8944 17196
rect 2372 17156 8944 17184
rect 2372 17144 2378 17156
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 20622 17184 20628 17196
rect 9088 17156 20628 17184
rect 9088 17144 9094 17156
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 25038 17144 25044 17196
rect 25096 17184 25102 17196
rect 43806 17184 43812 17196
rect 25096 17156 43812 17184
rect 25096 17144 25102 17156
rect 43806 17144 43812 17156
rect 43864 17144 43870 17196
rect 47762 17144 47768 17196
rect 47820 17184 47826 17196
rect 49694 17184 49700 17196
rect 47820 17156 49700 17184
rect 47820 17144 47826 17156
rect 49694 17144 49700 17156
rect 49752 17144 49758 17196
rect 49786 17144 49792 17196
rect 49844 17184 49850 17196
rect 55186 17184 55214 17224
rect 59998 17212 60004 17224
rect 60056 17212 60062 17264
rect 103698 17252 103704 17264
rect 65536 17224 103704 17252
rect 49844 17156 55214 17184
rect 49844 17144 49850 17156
rect 60826 17144 60832 17196
rect 60884 17184 60890 17196
rect 65536 17184 65564 17224
rect 103698 17212 103704 17224
rect 103756 17212 103762 17264
rect 104158 17212 104164 17264
rect 104216 17252 104222 17264
rect 111518 17252 111524 17264
rect 104216 17224 111524 17252
rect 104216 17212 104222 17224
rect 111518 17212 111524 17224
rect 111576 17212 111582 17264
rect 118878 17212 118884 17264
rect 118936 17252 118942 17264
rect 118936 17224 120810 17252
rect 118936 17212 118942 17224
rect 60884 17156 65564 17184
rect 60884 17144 60890 17156
rect 65886 17144 65892 17196
rect 65944 17184 65950 17196
rect 72142 17184 72148 17196
rect 65944 17156 72148 17184
rect 65944 17144 65950 17156
rect 72142 17144 72148 17156
rect 72200 17144 72206 17196
rect 78122 17144 78128 17196
rect 78180 17184 78186 17196
rect 82354 17184 82360 17196
rect 78180 17156 82360 17184
rect 78180 17144 78186 17156
rect 82354 17144 82360 17156
rect 82412 17144 82418 17196
rect 88794 17144 88800 17196
rect 88852 17184 88858 17196
rect 91370 17184 91376 17196
rect 88852 17156 91376 17184
rect 88852 17144 88858 17156
rect 91370 17144 91376 17156
rect 91428 17144 91434 17196
rect 95050 17144 95056 17196
rect 95108 17184 95114 17196
rect 101490 17184 101496 17196
rect 95108 17156 101496 17184
rect 95108 17144 95114 17156
rect 101490 17144 101496 17156
rect 101548 17144 101554 17196
rect 114554 17184 114560 17196
rect 103486 17156 114560 17184
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 26234 17116 26240 17128
rect 10836 17088 26240 17116
rect 10836 17076 10842 17088
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 42058 17076 42064 17128
rect 42116 17116 42122 17128
rect 46014 17116 46020 17128
rect 42116 17088 46020 17116
rect 42116 17076 42122 17088
rect 46014 17076 46020 17088
rect 46072 17076 46078 17128
rect 48866 17076 48872 17128
rect 48924 17116 48930 17128
rect 54570 17116 54576 17128
rect 48924 17088 54576 17116
rect 48924 17076 48930 17088
rect 54570 17076 54576 17088
rect 54628 17076 54634 17128
rect 56502 17076 56508 17128
rect 56560 17116 56566 17128
rect 65518 17116 65524 17128
rect 56560 17088 65524 17116
rect 56560 17076 56566 17088
rect 65518 17076 65524 17088
rect 65576 17076 65582 17128
rect 65702 17076 65708 17128
rect 65760 17116 65766 17128
rect 73982 17116 73988 17128
rect 65760 17088 73988 17116
rect 65760 17076 65766 17088
rect 73982 17076 73988 17088
rect 74040 17076 74046 17128
rect 88242 17076 88248 17128
rect 88300 17116 88306 17128
rect 93762 17116 93768 17128
rect 88300 17088 93768 17116
rect 88300 17076 88306 17088
rect 93762 17076 93768 17088
rect 93820 17076 93826 17128
rect 95694 17076 95700 17128
rect 95752 17116 95758 17128
rect 103486 17116 103514 17156
rect 114554 17144 114560 17156
rect 114612 17144 114618 17196
rect 120782 17184 120810 17224
rect 120902 17212 120908 17264
rect 120960 17252 120966 17264
rect 471974 17252 471980 17264
rect 120960 17224 471980 17252
rect 120960 17212 120966 17224
rect 471974 17212 471980 17224
rect 472032 17212 472038 17264
rect 126882 17184 126888 17196
rect 120782 17156 126888 17184
rect 126882 17144 126888 17156
rect 126940 17144 126946 17196
rect 142154 17184 142160 17196
rect 132466 17156 142160 17184
rect 95752 17088 103514 17116
rect 95752 17076 95758 17088
rect 104526 17076 104532 17128
rect 104584 17116 104590 17128
rect 114002 17116 114008 17128
rect 104584 17088 114008 17116
rect 104584 17076 104590 17088
rect 114002 17076 114008 17088
rect 114060 17076 114066 17128
rect 121730 17076 121736 17128
rect 121788 17116 121794 17128
rect 132466 17116 132494 17156
rect 142154 17144 142160 17156
rect 142212 17144 142218 17196
rect 143626 17144 143632 17196
rect 143684 17184 143690 17196
rect 151538 17184 151544 17196
rect 143684 17156 151544 17184
rect 143684 17144 143690 17156
rect 151538 17144 151544 17156
rect 151596 17144 151602 17196
rect 160186 17144 160192 17196
rect 160244 17184 160250 17196
rect 233510 17184 233516 17196
rect 160244 17156 233516 17184
rect 160244 17144 160250 17156
rect 233510 17144 233516 17156
rect 233568 17144 233574 17196
rect 121788 17088 132494 17116
rect 121788 17076 121794 17088
rect 476758 17076 476764 17128
rect 476816 17116 476822 17128
rect 480254 17116 480260 17128
rect 476816 17088 480260 17116
rect 476816 17076 476822 17088
rect 480254 17076 480260 17088
rect 480312 17076 480318 17128
rect 7742 17008 7748 17060
rect 7800 17048 7806 17060
rect 18414 17048 18420 17060
rect 7800 17020 18420 17048
rect 7800 17008 7806 17020
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 42150 17008 42156 17060
rect 42208 17048 42214 17060
rect 45830 17048 45836 17060
rect 42208 17020 45836 17048
rect 42208 17008 42214 17020
rect 45830 17008 45836 17020
rect 45888 17008 45894 17060
rect 48130 17008 48136 17060
rect 48188 17048 48194 17060
rect 50522 17048 50528 17060
rect 48188 17020 50528 17048
rect 48188 17008 48194 17020
rect 50522 17008 50528 17020
rect 50580 17008 50586 17060
rect 53650 17008 53656 17060
rect 53708 17048 53714 17060
rect 54938 17048 54944 17060
rect 53708 17020 54944 17048
rect 53708 17008 53714 17020
rect 54938 17008 54944 17020
rect 54996 17008 55002 17060
rect 71866 17008 71872 17060
rect 71924 17048 71930 17060
rect 95142 17048 95148 17060
rect 71924 17020 95148 17048
rect 71924 17008 71930 17020
rect 95142 17008 95148 17020
rect 95200 17008 95206 17060
rect 102318 17008 102324 17060
rect 102376 17048 102382 17060
rect 108298 17048 108304 17060
rect 102376 17020 108304 17048
rect 102376 17008 102382 17020
rect 108298 17008 108304 17020
rect 108356 17008 108362 17060
rect 110782 17008 110788 17060
rect 110840 17048 110846 17060
rect 117682 17048 117688 17060
rect 110840 17020 117688 17048
rect 110840 17008 110846 17020
rect 117682 17008 117688 17020
rect 117740 17008 117746 17060
rect 126146 17008 126152 17060
rect 126204 17048 126210 17060
rect 131114 17048 131120 17060
rect 126204 17020 131120 17048
rect 126204 17008 126210 17020
rect 131114 17008 131120 17020
rect 131172 17008 131178 17060
rect 146294 17008 146300 17060
rect 146352 17048 146358 17060
rect 149146 17048 149152 17060
rect 146352 17020 149152 17048
rect 146352 17008 146358 17020
rect 149146 17008 149152 17020
rect 149204 17008 149210 17060
rect 417510 17008 417516 17060
rect 417568 17048 417574 17060
rect 423674 17048 423680 17060
rect 417568 17020 423680 17048
rect 417568 17008 417574 17020
rect 423674 17008 423680 17020
rect 423732 17008 423738 17060
rect 438854 17008 438860 17060
rect 438912 17048 438918 17060
rect 441982 17048 441988 17060
rect 438912 17020 441988 17048
rect 438912 17008 438918 17020
rect 441982 17008 441988 17020
rect 442040 17008 442046 17060
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 40862 16980 40868 16992
rect 6052 16952 40868 16980
rect 6052 16940 6058 16952
rect 40862 16940 40868 16952
rect 40920 16940 40926 16992
rect 44174 16940 44180 16992
rect 44232 16980 44238 16992
rect 46750 16980 46756 16992
rect 44232 16952 46756 16980
rect 44232 16940 44238 16952
rect 46750 16940 46756 16952
rect 46808 16940 46814 16992
rect 48682 16940 48688 16992
rect 48740 16980 48746 16992
rect 54754 16980 54760 16992
rect 48740 16952 54760 16980
rect 48740 16940 48746 16952
rect 54754 16940 54760 16952
rect 54812 16940 54818 16992
rect 64138 16940 64144 16992
rect 64196 16980 64202 16992
rect 82814 16980 82820 16992
rect 64196 16952 82820 16980
rect 64196 16940 64202 16952
rect 82814 16940 82820 16952
rect 82872 16940 82878 16992
rect 83826 16940 83832 16992
rect 83884 16980 83890 16992
rect 84838 16980 84844 16992
rect 83884 16952 84844 16980
rect 83884 16940 83890 16952
rect 84838 16940 84844 16952
rect 84896 16940 84902 16992
rect 91002 16940 91008 16992
rect 91060 16980 91066 16992
rect 97810 16980 97816 16992
rect 91060 16952 97816 16980
rect 91060 16940 91066 16952
rect 97810 16940 97816 16952
rect 97868 16940 97874 16992
rect 100754 16940 100760 16992
rect 100812 16980 100818 16992
rect 112990 16980 112996 16992
rect 100812 16952 112996 16980
rect 100812 16940 100818 16952
rect 112990 16940 112996 16952
rect 113048 16940 113054 16992
rect 114462 16940 114468 16992
rect 114520 16980 114526 16992
rect 122374 16980 122380 16992
rect 114520 16952 122380 16980
rect 114520 16940 114526 16952
rect 122374 16940 122380 16952
rect 122432 16940 122438 16992
rect 17770 16872 17776 16924
rect 17828 16912 17834 16924
rect 72694 16912 72700 16924
rect 17828 16884 72700 16912
rect 17828 16872 17834 16884
rect 72694 16872 72700 16884
rect 72752 16872 72758 16924
rect 73338 16872 73344 16924
rect 73396 16912 73402 16924
rect 85482 16912 85488 16924
rect 73396 16884 85488 16912
rect 73396 16872 73402 16884
rect 85482 16872 85488 16884
rect 85540 16872 85546 16924
rect 91186 16872 91192 16924
rect 91244 16912 91250 16924
rect 93578 16912 93584 16924
rect 91244 16884 93584 16912
rect 91244 16872 91250 16884
rect 93578 16872 93584 16884
rect 93636 16872 93642 16924
rect 93762 16872 93768 16924
rect 93820 16912 93826 16924
rect 106090 16912 106096 16924
rect 93820 16884 106096 16912
rect 93820 16872 93826 16884
rect 106090 16872 106096 16884
rect 106148 16872 106154 16924
rect 113450 16872 113456 16924
rect 113508 16912 113514 16924
rect 120902 16912 120908 16924
rect 113508 16884 120908 16912
rect 113508 16872 113514 16884
rect 120902 16872 120908 16884
rect 120960 16872 120966 16924
rect 20070 16804 20076 16856
rect 20128 16844 20134 16856
rect 27614 16844 27620 16856
rect 20128 16816 27620 16844
rect 20128 16804 20134 16816
rect 27614 16804 27620 16816
rect 27672 16804 27678 16856
rect 43530 16804 43536 16856
rect 43588 16844 43594 16856
rect 45646 16844 45652 16856
rect 43588 16816 45652 16844
rect 43588 16804 43594 16816
rect 45646 16804 45652 16816
rect 45704 16804 45710 16856
rect 51442 16804 51448 16856
rect 51500 16844 51506 16856
rect 56042 16844 56048 16856
rect 51500 16816 56048 16844
rect 51500 16804 51506 16816
rect 56042 16804 56048 16816
rect 56100 16804 56106 16856
rect 67818 16804 67824 16856
rect 67876 16844 67882 16856
rect 70118 16844 70124 16856
rect 67876 16816 70124 16844
rect 67876 16804 67882 16816
rect 70118 16804 70124 16816
rect 70176 16804 70182 16856
rect 85850 16804 85856 16856
rect 85908 16844 85914 16856
rect 91002 16844 91008 16856
rect 85908 16816 91008 16844
rect 85908 16804 85914 16816
rect 91002 16804 91008 16816
rect 91060 16804 91066 16856
rect 91738 16804 91744 16856
rect 91796 16844 91802 16856
rect 96706 16844 96712 16856
rect 91796 16816 96712 16844
rect 91796 16804 91802 16816
rect 96706 16804 96712 16816
rect 96764 16804 96770 16856
rect 97810 16804 97816 16856
rect 97868 16844 97874 16856
rect 101306 16844 101312 16856
rect 97868 16816 101312 16844
rect 97868 16804 97874 16816
rect 101306 16804 101312 16816
rect 101364 16804 101370 16856
rect 102410 16804 102416 16856
rect 102468 16844 102474 16856
rect 106918 16844 106924 16856
rect 102468 16816 106924 16844
rect 102468 16804 102474 16816
rect 106918 16804 106924 16816
rect 106976 16804 106982 16856
rect 115106 16804 115112 16856
rect 115164 16844 115170 16856
rect 117498 16844 117504 16856
rect 115164 16816 117504 16844
rect 115164 16804 115170 16816
rect 117498 16804 117504 16816
rect 117556 16804 117562 16856
rect 437474 16804 437480 16856
rect 437532 16844 437538 16856
rect 441614 16844 441620 16856
rect 437532 16816 441620 16844
rect 437532 16804 437538 16816
rect 441614 16804 441620 16816
rect 441672 16804 441678 16856
rect 43622 16736 43628 16788
rect 43680 16776 43686 16788
rect 46198 16776 46204 16788
rect 43680 16748 46204 16776
rect 43680 16736 43686 16748
rect 46198 16736 46204 16748
rect 46256 16736 46262 16788
rect 52546 16736 52552 16788
rect 52604 16776 52610 16788
rect 55858 16776 55864 16788
rect 52604 16748 55864 16776
rect 52604 16736 52610 16748
rect 55858 16736 55864 16748
rect 55916 16736 55922 16788
rect 66438 16736 66444 16788
rect 66496 16776 66502 16788
rect 67910 16776 67916 16788
rect 66496 16748 67916 16776
rect 66496 16736 66502 16748
rect 67910 16736 67916 16748
rect 67968 16736 67974 16788
rect 81618 16736 81624 16788
rect 81676 16776 81682 16788
rect 84470 16776 84476 16788
rect 81676 16748 84476 16776
rect 81676 16736 81682 16748
rect 84470 16736 84476 16748
rect 84528 16736 84534 16788
rect 111242 16736 111248 16788
rect 111300 16776 111306 16788
rect 242802 16776 242808 16788
rect 111300 16748 242808 16776
rect 111300 16736 111306 16748
rect 242802 16736 242808 16748
rect 242860 16736 242866 16788
rect 39298 16668 39304 16720
rect 39356 16708 39362 16720
rect 45462 16708 45468 16720
rect 39356 16680 45468 16708
rect 39356 16668 39362 16680
rect 45462 16668 45468 16680
rect 45520 16668 45526 16720
rect 61654 16668 61660 16720
rect 61712 16708 61718 16720
rect 66806 16708 66812 16720
rect 61712 16680 66812 16708
rect 61712 16668 61718 16680
rect 66806 16668 66812 16680
rect 66864 16668 66870 16720
rect 71774 16668 71780 16720
rect 71832 16708 71838 16720
rect 71832 16680 79364 16708
rect 71832 16668 71838 16680
rect 934 16600 940 16652
rect 992 16640 998 16652
rect 8386 16640 8392 16652
rect 992 16612 8392 16640
rect 992 16600 998 16612
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 44818 16600 44824 16652
rect 44876 16640 44882 16652
rect 46382 16640 46388 16652
rect 44876 16612 46388 16640
rect 44876 16600 44882 16612
rect 46382 16600 46388 16612
rect 46440 16600 46446 16652
rect 61746 16600 61752 16652
rect 61804 16640 61810 16652
rect 64138 16640 64144 16652
rect 61804 16612 64144 16640
rect 61804 16600 61810 16612
rect 64138 16600 64144 16612
rect 64196 16600 64202 16652
rect 64506 16600 64512 16652
rect 64564 16640 64570 16652
rect 65610 16640 65616 16652
rect 64564 16612 65616 16640
rect 64564 16600 64570 16612
rect 65610 16600 65616 16612
rect 65668 16600 65674 16652
rect 66346 16600 66352 16652
rect 66404 16640 66410 16652
rect 68278 16640 68284 16652
rect 66404 16612 68284 16640
rect 66404 16600 66410 16612
rect 68278 16600 68284 16612
rect 68336 16600 68342 16652
rect 72418 16600 72424 16652
rect 72476 16640 72482 16652
rect 76742 16640 76748 16652
rect 72476 16612 76748 16640
rect 72476 16600 72482 16612
rect 76742 16600 76748 16612
rect 76800 16600 76806 16652
rect 79336 16640 79364 16680
rect 82906 16668 82912 16720
rect 82964 16708 82970 16720
rect 85114 16708 85120 16720
rect 82964 16680 85120 16708
rect 82964 16668 82970 16680
rect 85114 16668 85120 16680
rect 85172 16668 85178 16720
rect 93394 16668 93400 16720
rect 93452 16708 93458 16720
rect 94682 16708 94688 16720
rect 93452 16680 94688 16708
rect 93452 16668 93458 16680
rect 94682 16668 94688 16680
rect 94740 16668 94746 16720
rect 97626 16668 97632 16720
rect 97684 16708 97690 16720
rect 104618 16708 104624 16720
rect 97684 16680 104624 16708
rect 97684 16668 97690 16680
rect 104618 16668 104624 16680
rect 104676 16668 104682 16720
rect 107930 16668 107936 16720
rect 107988 16708 107994 16720
rect 240226 16708 240232 16720
rect 107988 16680 240232 16708
rect 107988 16668 107994 16680
rect 240226 16668 240232 16680
rect 240284 16668 240290 16720
rect 97902 16640 97908 16652
rect 79336 16612 97908 16640
rect 97902 16600 97908 16612
rect 97960 16600 97966 16652
rect 116118 16600 116124 16652
rect 116176 16640 116182 16652
rect 116176 16612 118694 16640
rect 116176 16600 116182 16612
rect 7926 16532 7932 16584
rect 7984 16572 7990 16584
rect 11054 16572 11060 16584
rect 7984 16544 11060 16572
rect 7984 16532 7990 16544
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 70486 16572 70492 16584
rect 12406 16544 70492 16572
rect 10870 16464 10876 16516
rect 10928 16504 10934 16516
rect 12406 16504 12434 16544
rect 70486 16532 70492 16544
rect 70544 16532 70550 16584
rect 116394 16532 116400 16584
rect 116452 16572 116458 16584
rect 116854 16572 116860 16584
rect 116452 16544 116860 16572
rect 116452 16532 116458 16544
rect 116854 16532 116860 16544
rect 116912 16532 116918 16584
rect 118666 16572 118694 16612
rect 122650 16600 122656 16652
rect 122708 16640 122714 16652
rect 123754 16640 123760 16652
rect 122708 16612 123760 16640
rect 122708 16600 122714 16612
rect 123754 16600 123760 16612
rect 123812 16600 123818 16652
rect 129734 16600 129740 16652
rect 129792 16640 129798 16652
rect 132494 16640 132500 16652
rect 129792 16612 132500 16640
rect 129792 16600 129798 16612
rect 132494 16600 132500 16612
rect 132552 16600 132558 16652
rect 153654 16600 153660 16652
rect 153712 16640 153718 16652
rect 153930 16640 153936 16652
rect 153712 16612 153936 16640
rect 153712 16600 153718 16612
rect 153930 16600 153936 16612
rect 153988 16600 153994 16652
rect 121178 16572 121184 16584
rect 118666 16544 121184 16572
rect 121178 16532 121184 16544
rect 121236 16532 121242 16584
rect 129550 16532 129556 16584
rect 129608 16572 129614 16584
rect 133782 16572 133788 16584
rect 129608 16544 133788 16572
rect 129608 16532 129614 16544
rect 133782 16532 133788 16544
rect 133840 16532 133846 16584
rect 142154 16532 142160 16584
rect 142212 16572 142218 16584
rect 147674 16572 147680 16584
rect 142212 16544 147680 16572
rect 142212 16532 142218 16544
rect 147674 16532 147680 16544
rect 147732 16532 147738 16584
rect 158254 16572 158260 16584
rect 151786 16544 158260 16572
rect 10928 16476 12434 16504
rect 10928 16464 10934 16476
rect 16482 16464 16488 16516
rect 16540 16504 16546 16516
rect 18966 16504 18972 16516
rect 16540 16476 18972 16504
rect 16540 16464 16546 16476
rect 18966 16464 18972 16476
rect 19024 16464 19030 16516
rect 66254 16504 66260 16516
rect 21376 16476 66260 16504
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 21376 16436 21404 16476
rect 66254 16464 66260 16476
rect 66312 16464 66318 16516
rect 83918 16464 83924 16516
rect 83976 16504 83982 16516
rect 86494 16504 86500 16516
rect 83976 16476 86500 16504
rect 83976 16464 83982 16476
rect 86494 16464 86500 16476
rect 86552 16464 86558 16516
rect 111058 16464 111064 16516
rect 111116 16504 111122 16516
rect 117314 16504 117320 16516
rect 111116 16476 117320 16504
rect 111116 16464 111122 16476
rect 117314 16464 117320 16476
rect 117372 16464 117378 16516
rect 143534 16464 143540 16516
rect 143592 16504 143598 16516
rect 151786 16504 151814 16544
rect 158254 16532 158260 16544
rect 158312 16532 158318 16584
rect 143592 16476 151814 16504
rect 143592 16464 143598 16476
rect 10652 16408 21404 16436
rect 10652 16396 10658 16408
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 96890 16436 96896 16448
rect 26292 16408 96896 16436
rect 26292 16396 26298 16408
rect 96890 16396 96896 16408
rect 96948 16396 96954 16448
rect 99282 16396 99288 16448
rect 99340 16436 99346 16448
rect 201402 16436 201408 16448
rect 99340 16408 201408 16436
rect 99340 16396 99346 16408
rect 201402 16396 201408 16408
rect 201460 16396 201466 16448
rect 212810 16396 212816 16448
rect 212868 16436 212874 16448
rect 295334 16436 295340 16448
rect 212868 16408 295340 16436
rect 212868 16396 212874 16408
rect 295334 16396 295340 16408
rect 295392 16396 295398 16448
rect 6730 16328 6736 16380
rect 6788 16368 6794 16380
rect 15470 16368 15476 16380
rect 6788 16340 15476 16368
rect 6788 16328 6794 16340
rect 15470 16328 15476 16340
rect 15528 16328 15534 16380
rect 24854 16328 24860 16380
rect 24912 16368 24918 16380
rect 91738 16368 91744 16380
rect 24912 16340 91744 16368
rect 24912 16328 24918 16340
rect 91738 16328 91744 16340
rect 91796 16328 91802 16380
rect 95510 16328 95516 16380
rect 95568 16368 95574 16380
rect 262490 16368 262496 16380
rect 95568 16340 262496 16368
rect 95568 16328 95574 16340
rect 262490 16328 262496 16340
rect 262548 16328 262554 16380
rect 267826 16328 267832 16380
rect 267884 16368 267890 16380
rect 280338 16368 280344 16380
rect 267884 16340 280344 16368
rect 267884 16328 267890 16340
rect 280338 16328 280344 16340
rect 280396 16328 280402 16380
rect 280430 16328 280436 16380
rect 280488 16368 280494 16380
rect 380894 16368 380900 16380
rect 280488 16340 380900 16368
rect 280488 16328 280494 16340
rect 380894 16328 380900 16340
rect 380952 16328 380958 16380
rect 6454 16260 6460 16312
rect 6512 16300 6518 16312
rect 19242 16300 19248 16312
rect 6512 16272 19248 16300
rect 6512 16260 6518 16272
rect 19242 16260 19248 16272
rect 19300 16260 19306 16312
rect 21358 16260 21364 16312
rect 21416 16300 21422 16312
rect 71038 16300 71044 16312
rect 21416 16272 71044 16300
rect 21416 16260 21422 16272
rect 71038 16260 71044 16272
rect 71096 16260 71102 16312
rect 71866 16260 71872 16312
rect 71924 16300 71930 16312
rect 79502 16300 79508 16312
rect 71924 16272 79508 16300
rect 71924 16260 71930 16272
rect 79502 16260 79508 16272
rect 79560 16260 79566 16312
rect 112898 16260 112904 16312
rect 112956 16300 112962 16312
rect 117222 16300 117228 16312
rect 112956 16272 117228 16300
rect 112956 16260 112962 16272
rect 117222 16260 117228 16272
rect 117280 16260 117286 16312
rect 117314 16260 117320 16312
rect 117372 16300 117378 16312
rect 291746 16300 291752 16312
rect 117372 16272 291752 16300
rect 117372 16260 117378 16272
rect 291746 16260 291752 16272
rect 291804 16260 291810 16312
rect 391290 16260 391296 16312
rect 391348 16300 391354 16312
rect 399018 16300 399024 16312
rect 391348 16272 399024 16300
rect 391348 16260 391354 16272
rect 399018 16260 399024 16272
rect 399076 16260 399082 16312
rect 15194 16192 15200 16244
rect 15252 16232 15258 16244
rect 43346 16232 43352 16244
rect 15252 16204 43352 16232
rect 15252 16192 15258 16204
rect 43346 16192 43352 16204
rect 43404 16192 43410 16244
rect 55582 16192 55588 16244
rect 55640 16232 55646 16244
rect 73798 16232 73804 16244
rect 55640 16204 73804 16232
rect 55640 16192 55646 16204
rect 73798 16192 73804 16204
rect 73856 16192 73862 16244
rect 90818 16192 90824 16244
rect 90876 16232 90882 16244
rect 283006 16232 283012 16244
rect 90876 16204 283012 16232
rect 90876 16192 90882 16204
rect 283006 16192 283012 16204
rect 283064 16192 283070 16244
rect 294598 16192 294604 16244
rect 294656 16232 294662 16244
rect 417326 16232 417332 16244
rect 294656 16204 417332 16232
rect 294656 16192 294662 16204
rect 417326 16192 417332 16204
rect 417384 16192 417390 16244
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 41598 16164 41604 16176
rect 13136 16136 41604 16164
rect 13136 16124 13142 16136
rect 41598 16124 41604 16136
rect 41656 16124 41662 16176
rect 47302 16124 47308 16176
rect 47360 16164 47366 16176
rect 74534 16164 74540 16176
rect 47360 16136 74540 16164
rect 47360 16124 47366 16136
rect 74534 16124 74540 16136
rect 74592 16124 74598 16176
rect 77018 16124 77024 16176
rect 77076 16164 77082 16176
rect 81526 16164 81532 16176
rect 77076 16136 81532 16164
rect 77076 16124 77082 16136
rect 81526 16124 81532 16136
rect 81584 16124 81590 16176
rect 82446 16124 82452 16176
rect 82504 16164 82510 16176
rect 87690 16164 87696 16176
rect 82504 16136 87696 16164
rect 82504 16124 82510 16136
rect 87690 16124 87696 16136
rect 87748 16124 87754 16176
rect 89438 16124 89444 16176
rect 89496 16164 89502 16176
rect 223482 16164 223488 16176
rect 89496 16136 223488 16164
rect 89496 16124 89502 16136
rect 223482 16124 223488 16136
rect 223540 16124 223546 16176
rect 240226 16124 240232 16176
rect 240284 16164 240290 16176
rect 436738 16164 436744 16176
rect 240284 16136 436744 16164
rect 240284 16124 240290 16136
rect 436738 16124 436744 16136
rect 436796 16124 436802 16176
rect 7650 16056 7656 16108
rect 7708 16096 7714 16108
rect 41046 16096 41052 16108
rect 7708 16068 41052 16096
rect 7708 16056 7714 16068
rect 41046 16056 41052 16068
rect 41104 16056 41110 16108
rect 53926 16056 53932 16108
rect 53984 16096 53990 16108
rect 86954 16096 86960 16108
rect 53984 16068 86960 16096
rect 53984 16056 53990 16068
rect 86954 16056 86960 16068
rect 87012 16056 87018 16108
rect 91278 16056 91284 16108
rect 91336 16096 91342 16108
rect 327718 16096 327724 16108
rect 91336 16068 327724 16096
rect 91336 16056 91342 16068
rect 327718 16056 327724 16068
rect 327776 16056 327782 16108
rect 372614 16056 372620 16108
rect 372672 16096 372678 16108
rect 377766 16096 377772 16108
rect 372672 16068 377772 16096
rect 372672 16056 372678 16068
rect 377766 16056 377772 16068
rect 377824 16056 377830 16108
rect 381538 16056 381544 16108
rect 381596 16096 381602 16108
rect 395798 16096 395804 16108
rect 381596 16068 395804 16096
rect 381596 16056 381602 16068
rect 395798 16056 395804 16068
rect 395856 16056 395862 16108
rect 399478 16056 399484 16108
rect 399536 16096 399542 16108
rect 438854 16096 438860 16108
rect 399536 16068 438860 16096
rect 399536 16056 399542 16068
rect 438854 16056 438860 16068
rect 438912 16056 438918 16108
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 39942 16028 39948 16040
rect 4856 16000 39948 16028
rect 4856 15988 4862 16000
rect 39942 15988 39948 16000
rect 40000 15988 40006 16040
rect 55398 15988 55404 16040
rect 55456 16028 55462 16040
rect 97258 16028 97264 16040
rect 55456 16000 97264 16028
rect 55456 15988 55462 16000
rect 97258 15988 97264 16000
rect 97316 15988 97322 16040
rect 98270 15988 98276 16040
rect 98328 16028 98334 16040
rect 374086 16028 374092 16040
rect 98328 16000 374092 16028
rect 98328 15988 98334 16000
rect 374086 15988 374092 16000
rect 374144 15988 374150 16040
rect 381906 15988 381912 16040
rect 381964 16028 381970 16040
rect 390646 16028 390652 16040
rect 381964 16000 390652 16028
rect 381964 15988 381970 16000
rect 390646 15988 390652 16000
rect 390704 15988 390710 16040
rect 395338 15988 395344 16040
rect 395396 16028 395402 16040
rect 476758 16028 476764 16040
rect 395396 16000 476764 16028
rect 395396 15988 395402 16000
rect 476758 15988 476764 16000
rect 476816 15988 476822 16040
rect 5166 15920 5172 15972
rect 5224 15960 5230 15972
rect 20898 15960 20904 15972
rect 5224 15932 20904 15960
rect 5224 15920 5230 15932
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 59170 15960 59176 15972
rect 23440 15932 59176 15960
rect 23440 15920 23446 15932
rect 59170 15920 59176 15932
rect 59228 15920 59234 15972
rect 63770 15920 63776 15972
rect 63828 15960 63834 15972
rect 66162 15960 66168 15972
rect 63828 15932 66168 15960
rect 63828 15920 63834 15932
rect 66162 15920 66168 15932
rect 66220 15920 66226 15972
rect 66254 15920 66260 15972
rect 66312 15960 66318 15972
rect 111886 15960 111892 15972
rect 66312 15932 111892 15960
rect 66312 15920 66318 15932
rect 111886 15920 111892 15932
rect 111944 15920 111950 15972
rect 114370 15920 114376 15972
rect 114428 15960 114434 15972
rect 478138 15960 478144 15972
rect 114428 15932 478144 15960
rect 114428 15920 114434 15932
rect 478138 15920 478144 15932
rect 478196 15920 478202 15972
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 40126 15892 40132 15904
rect 3476 15864 40132 15892
rect 3476 15852 3482 15864
rect 40126 15852 40132 15864
rect 40184 15852 40190 15904
rect 57606 15852 57612 15904
rect 57664 15892 57670 15904
rect 111058 15892 111064 15904
rect 57664 15864 111064 15892
rect 57664 15852 57670 15864
rect 111058 15852 111064 15864
rect 111116 15852 111122 15904
rect 116762 15852 116768 15904
rect 116820 15892 116826 15904
rect 485130 15892 485136 15904
rect 116820 15864 485136 15892
rect 116820 15852 116826 15864
rect 485130 15852 485136 15864
rect 485188 15852 485194 15904
rect 13722 15784 13728 15836
rect 13780 15824 13786 15836
rect 15746 15824 15752 15836
rect 13780 15796 15752 15824
rect 13780 15784 13786 15796
rect 15746 15784 15752 15796
rect 15804 15784 15810 15836
rect 17862 15784 17868 15836
rect 17920 15824 17926 15836
rect 33686 15824 33692 15836
rect 17920 15796 33692 15824
rect 17920 15784 17926 15796
rect 33686 15784 33692 15796
rect 33744 15784 33750 15836
rect 56318 15784 56324 15836
rect 56376 15824 56382 15836
rect 91738 15824 91744 15836
rect 56376 15796 91744 15824
rect 56376 15784 56382 15796
rect 91738 15784 91744 15796
rect 91796 15784 91802 15836
rect 92014 15784 92020 15836
rect 92072 15824 92078 15836
rect 98270 15824 98276 15836
rect 92072 15796 98276 15824
rect 92072 15784 92078 15796
rect 98270 15784 98276 15796
rect 98328 15784 98334 15836
rect 102962 15784 102968 15836
rect 103020 15824 103026 15836
rect 107562 15824 107568 15836
rect 103020 15796 107568 15824
rect 103020 15784 103026 15796
rect 107562 15784 107568 15796
rect 107620 15784 107626 15836
rect 109402 15784 109408 15836
rect 109460 15824 109466 15836
rect 143626 15824 143632 15836
rect 109460 15796 143632 15824
rect 109460 15784 109466 15796
rect 143626 15784 143632 15796
rect 143684 15784 143690 15836
rect 150434 15784 150440 15836
rect 150492 15824 150498 15836
rect 158162 15824 158168 15836
rect 150492 15796 158168 15824
rect 150492 15784 150498 15796
rect 158162 15784 158168 15796
rect 158220 15784 158226 15836
rect 13538 15716 13544 15768
rect 13596 15756 13602 15768
rect 22094 15756 22100 15768
rect 13596 15728 22100 15756
rect 13596 15716 13602 15728
rect 22094 15716 22100 15728
rect 22152 15716 22158 15768
rect 50062 15716 50068 15768
rect 50120 15756 50126 15768
rect 50120 15728 61976 15756
rect 50120 15716 50126 15728
rect 53190 15648 53196 15700
rect 53248 15688 53254 15700
rect 61562 15688 61568 15700
rect 53248 15660 61568 15688
rect 53248 15648 53254 15660
rect 61562 15648 61568 15660
rect 61620 15648 61626 15700
rect 61948 15688 61976 15728
rect 62022 15716 62028 15768
rect 62080 15756 62086 15768
rect 66254 15756 66260 15768
rect 62080 15728 66260 15756
rect 62080 15716 62086 15728
rect 66254 15716 66260 15728
rect 66312 15716 66318 15768
rect 73614 15716 73620 15768
rect 73672 15756 73678 15768
rect 81434 15756 81440 15768
rect 73672 15728 81440 15756
rect 73672 15716 73678 15728
rect 81434 15716 81440 15728
rect 81492 15716 81498 15768
rect 91002 15716 91008 15768
rect 91060 15756 91066 15768
rect 118142 15756 118148 15768
rect 91060 15728 118148 15756
rect 91060 15716 91066 15728
rect 118142 15716 118148 15728
rect 118200 15716 118206 15768
rect 122742 15716 122748 15768
rect 122800 15756 122806 15768
rect 123570 15756 123576 15768
rect 122800 15728 123576 15756
rect 122800 15716 122806 15728
rect 123570 15716 123576 15728
rect 123628 15716 123634 15768
rect 153102 15756 153108 15768
rect 127636 15728 153108 15756
rect 65058 15688 65064 15700
rect 61948 15660 65064 15688
rect 65058 15648 65064 15660
rect 65116 15648 65122 15700
rect 90358 15648 90364 15700
rect 90416 15688 90422 15700
rect 98086 15688 98092 15700
rect 90416 15660 98092 15688
rect 90416 15648 90422 15660
rect 98086 15648 98092 15660
rect 98144 15648 98150 15700
rect 99190 15648 99196 15700
rect 99248 15688 99254 15700
rect 112530 15688 112536 15700
rect 99248 15660 112536 15688
rect 99248 15648 99254 15660
rect 112530 15648 112536 15660
rect 112588 15648 112594 15700
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 20530 15620 20536 15632
rect 15436 15592 20536 15620
rect 15436 15580 15442 15592
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 84102 15580 84108 15632
rect 84160 15620 84166 15632
rect 89898 15620 89904 15632
rect 84160 15592 89904 15620
rect 84160 15580 84166 15592
rect 89898 15580 89904 15592
rect 89956 15580 89962 15632
rect 97718 15580 97724 15632
rect 97776 15620 97782 15632
rect 98178 15620 98184 15632
rect 97776 15592 98184 15620
rect 97776 15580 97782 15592
rect 98178 15580 98184 15592
rect 98236 15580 98242 15632
rect 18506 15512 18512 15564
rect 18564 15552 18570 15564
rect 22370 15552 22376 15564
rect 18564 15524 22376 15552
rect 18564 15512 18570 15524
rect 22370 15512 22376 15524
rect 22428 15512 22434 15564
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 45738 15484 45744 15496
rect 19668 15456 45744 15484
rect 19668 15444 19674 15456
rect 45738 15444 45744 15456
rect 45796 15444 45802 15496
rect 81710 15444 81716 15496
rect 81768 15484 81774 15496
rect 127636 15484 127664 15728
rect 153102 15716 153108 15728
rect 153160 15716 153166 15768
rect 132494 15648 132500 15700
rect 132552 15688 132558 15700
rect 143074 15688 143080 15700
rect 132552 15660 143080 15688
rect 132552 15648 132558 15660
rect 143074 15648 143080 15660
rect 143132 15648 143138 15700
rect 81768 15456 127664 15484
rect 81768 15444 81774 15456
rect 77846 15376 77852 15428
rect 77904 15416 77910 15428
rect 151998 15416 152004 15428
rect 77904 15388 152004 15416
rect 77904 15376 77910 15388
rect 151998 15376 152004 15388
rect 152056 15376 152062 15428
rect 65978 15308 65984 15360
rect 66036 15348 66042 15360
rect 167178 15348 167184 15360
rect 66036 15320 167184 15348
rect 66036 15308 66042 15320
rect 167178 15308 167184 15320
rect 167236 15308 167242 15360
rect 377582 15308 377588 15360
rect 377640 15348 377646 15360
rect 381170 15348 381176 15360
rect 377640 15320 381176 15348
rect 377640 15308 377646 15320
rect 381170 15308 381176 15320
rect 381228 15308 381234 15360
rect 18046 15240 18052 15292
rect 18104 15280 18110 15292
rect 20162 15280 20168 15292
rect 18104 15252 20168 15280
rect 18104 15240 18110 15252
rect 20162 15240 20168 15252
rect 20220 15240 20226 15292
rect 66070 15240 66076 15292
rect 66128 15280 66134 15292
rect 70486 15280 70492 15292
rect 66128 15252 70492 15280
rect 66128 15240 66134 15252
rect 70486 15240 70492 15252
rect 70544 15240 70550 15292
rect 86954 15240 86960 15292
rect 87012 15280 87018 15292
rect 89622 15280 89628 15292
rect 87012 15252 89628 15280
rect 87012 15240 87018 15252
rect 89622 15240 89628 15252
rect 89680 15240 89686 15292
rect 153102 15240 153108 15292
rect 153160 15280 153166 15292
rect 179506 15280 179512 15292
rect 153160 15252 179512 15280
rect 153160 15240 153166 15252
rect 179506 15240 179512 15252
rect 179564 15240 179570 15292
rect 16758 15172 16764 15224
rect 16816 15212 16822 15224
rect 24854 15212 24860 15224
rect 16816 15184 24860 15212
rect 16816 15172 16822 15184
rect 24854 15172 24860 15184
rect 24912 15172 24918 15224
rect 42242 15172 42248 15224
rect 42300 15212 42306 15224
rect 42886 15212 42892 15224
rect 42300 15184 42892 15212
rect 42300 15172 42306 15184
rect 42886 15172 42892 15184
rect 42944 15172 42950 15224
rect 60182 15172 60188 15224
rect 60240 15212 60246 15224
rect 61838 15212 61844 15224
rect 60240 15184 61844 15212
rect 60240 15172 60246 15184
rect 61838 15172 61844 15184
rect 61896 15172 61902 15224
rect 75638 15172 75644 15224
rect 75696 15212 75702 15224
rect 78490 15212 78496 15224
rect 75696 15184 78496 15212
rect 75696 15172 75702 15184
rect 78490 15172 78496 15184
rect 78548 15172 78554 15224
rect 81342 15172 81348 15224
rect 81400 15212 81406 15224
rect 82538 15212 82544 15224
rect 81400 15184 82544 15212
rect 81400 15172 81406 15184
rect 82538 15172 82544 15184
rect 82596 15172 82602 15224
rect 87782 15172 87788 15224
rect 87840 15212 87846 15224
rect 88978 15212 88984 15224
rect 87840 15184 88984 15212
rect 87840 15172 87846 15184
rect 88978 15172 88984 15184
rect 89036 15172 89042 15224
rect 90174 15172 90180 15224
rect 90232 15212 90238 15224
rect 92566 15212 92572 15224
rect 90232 15184 92572 15212
rect 90232 15172 90238 15184
rect 92566 15172 92572 15184
rect 92624 15172 92630 15224
rect 92750 15172 92756 15224
rect 92808 15212 92814 15224
rect 95786 15212 95792 15224
rect 92808 15184 95792 15212
rect 92808 15172 92814 15184
rect 95786 15172 95792 15184
rect 95844 15172 95850 15224
rect 99374 15172 99380 15224
rect 99432 15212 99438 15224
rect 101582 15212 101588 15224
rect 99432 15184 101588 15212
rect 99432 15172 99438 15184
rect 101582 15172 101588 15184
rect 101640 15172 101646 15224
rect 124306 15172 124312 15224
rect 124364 15212 124370 15224
rect 128538 15212 128544 15224
rect 124364 15184 128544 15212
rect 124364 15172 124370 15184
rect 128538 15172 128544 15184
rect 128596 15172 128602 15224
rect 130010 15172 130016 15224
rect 130068 15212 130074 15224
rect 130068 15184 132494 15212
rect 130068 15172 130074 15184
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 10778 15144 10784 15156
rect 4120 15116 10784 15144
rect 4120 15104 4126 15116
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 77294 15144 77300 15156
rect 13412 15116 77300 15144
rect 13412 15104 13418 15116
rect 77294 15104 77300 15116
rect 77352 15104 77358 15156
rect 122282 15104 122288 15156
rect 122340 15144 122346 15156
rect 124122 15144 124128 15156
rect 122340 15116 124128 15144
rect 122340 15104 122346 15116
rect 124122 15104 124128 15116
rect 124180 15104 124186 15156
rect 132466 15144 132494 15184
rect 155402 15172 155408 15224
rect 155460 15212 155466 15224
rect 532050 15212 532056 15224
rect 155460 15184 532056 15212
rect 155460 15172 155466 15184
rect 532050 15172 532056 15184
rect 532108 15172 532114 15224
rect 158438 15144 158444 15156
rect 132466 15116 158444 15144
rect 158438 15104 158444 15116
rect 158496 15104 158502 15156
rect 187602 15104 187608 15156
rect 187660 15144 187666 15156
rect 205082 15144 205088 15156
rect 187660 15116 205088 15144
rect 187660 15104 187666 15116
rect 205082 15104 205088 15116
rect 205140 15104 205146 15156
rect 8110 15036 8116 15088
rect 8168 15076 8174 15088
rect 15378 15076 15384 15088
rect 8168 15048 15384 15076
rect 8168 15036 8174 15048
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 64230 15076 64236 15088
rect 15488 15048 64236 15076
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 10594 15008 10600 15020
rect 2648 14980 10600 15008
rect 2648 14968 2654 14980
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 10962 14968 10968 15020
rect 11020 15008 11026 15020
rect 15488 15008 15516 15048
rect 64230 15036 64236 15048
rect 64288 15036 64294 15088
rect 64322 15036 64328 15088
rect 64380 15076 64386 15088
rect 65518 15076 65524 15088
rect 64380 15048 65524 15076
rect 64380 15036 64386 15048
rect 65518 15036 65524 15048
rect 65576 15036 65582 15088
rect 142246 15036 142252 15088
rect 142304 15076 142310 15088
rect 150434 15076 150440 15088
rect 142304 15048 150440 15076
rect 142304 15036 142310 15048
rect 150434 15036 150440 15048
rect 150492 15036 150498 15088
rect 89714 15008 89720 15020
rect 11020 14980 15516 15008
rect 16546 14980 89720 15008
rect 11020 14968 11026 14980
rect 2498 14900 2504 14952
rect 2556 14940 2562 14952
rect 10870 14940 10876 14952
rect 2556 14912 10876 14940
rect 2556 14900 2562 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 16546 14940 16574 14980
rect 89714 14968 89720 14980
rect 89772 14968 89778 15020
rect 131114 14968 131120 15020
rect 131172 15008 131178 15020
rect 243538 15008 243544 15020
rect 131172 14980 243544 15008
rect 131172 14968 131178 14980
rect 243538 14968 243544 14980
rect 243596 14968 243602 15020
rect 15804 14912 16574 14940
rect 15804 14900 15810 14912
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 19150 14940 19156 14952
rect 18932 14912 19156 14940
rect 18932 14900 18938 14912
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 58158 14900 58164 14952
rect 58216 14940 58222 14952
rect 58216 14912 65610 14940
rect 58216 14900 58222 14912
rect 3694 14832 3700 14884
rect 3752 14872 3758 14884
rect 15286 14872 15292 14884
rect 3752 14844 15292 14872
rect 3752 14832 3758 14844
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 62758 14872 62764 14884
rect 15436 14844 62764 14872
rect 15436 14832 15442 14844
rect 62758 14832 62764 14844
rect 62816 14832 62822 14884
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 19150 14804 19156 14816
rect 3844 14776 19156 14804
rect 3844 14764 3850 14776
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 65150 14804 65156 14816
rect 20680 14776 65156 14804
rect 20680 14764 20686 14776
rect 65150 14764 65156 14776
rect 65208 14764 65214 14816
rect 19242 14696 19248 14748
rect 19300 14736 19306 14748
rect 61654 14736 61660 14748
rect 19300 14708 61660 14736
rect 19300 14696 19306 14708
rect 61654 14696 61660 14708
rect 61712 14696 61718 14748
rect 4890 14628 4896 14680
rect 4948 14668 4954 14680
rect 18598 14668 18604 14680
rect 4948 14640 18604 14668
rect 4948 14628 4954 14640
rect 18598 14628 18604 14640
rect 18656 14628 18662 14680
rect 19886 14628 19892 14680
rect 19944 14668 19950 14680
rect 60642 14668 60648 14680
rect 19944 14640 60648 14668
rect 19944 14628 19950 14640
rect 60642 14628 60648 14640
rect 60700 14628 60706 14680
rect 65582 14668 65610 14912
rect 90542 14900 90548 14952
rect 90600 14940 90606 14952
rect 210970 14940 210976 14952
rect 90600 14912 210976 14940
rect 90600 14900 90606 14912
rect 210970 14900 210976 14912
rect 211028 14900 211034 14952
rect 349798 14900 349804 14952
rect 349856 14940 349862 14952
rect 390554 14940 390560 14952
rect 349856 14912 390560 14940
rect 349856 14900 349862 14912
rect 390554 14900 390560 14912
rect 390612 14900 390618 14952
rect 439406 14900 439412 14952
rect 439464 14940 439470 14952
rect 442902 14940 442908 14952
rect 439464 14912 442908 14940
rect 439464 14900 439470 14912
rect 442902 14900 442908 14912
rect 442960 14900 442966 14952
rect 449158 14900 449164 14952
rect 449216 14940 449222 14952
rect 456058 14940 456064 14952
rect 449216 14912 456064 14940
rect 449216 14900 449222 14912
rect 456058 14900 456064 14912
rect 456116 14900 456122 14952
rect 71406 14832 71412 14884
rect 71464 14872 71470 14884
rect 197354 14872 197360 14884
rect 71464 14844 197360 14872
rect 71464 14832 71470 14844
rect 197354 14832 197360 14844
rect 197412 14832 197418 14884
rect 242802 14832 242808 14884
rect 242860 14872 242866 14884
rect 263594 14872 263600 14884
rect 242860 14844 263600 14872
rect 242860 14832 242866 14844
rect 263594 14832 263600 14844
rect 263652 14832 263658 14884
rect 291746 14832 291752 14884
rect 291804 14872 291810 14884
rect 353294 14872 353300 14884
rect 291804 14844 353300 14872
rect 291804 14832 291810 14844
rect 353294 14832 353300 14844
rect 353352 14832 353358 14884
rect 399570 14832 399576 14884
rect 399628 14872 399634 14884
rect 413554 14872 413560 14884
rect 399628 14844 413560 14872
rect 399628 14832 399634 14844
rect 413554 14832 413560 14844
rect 413612 14832 413618 14884
rect 477402 14832 477408 14884
rect 477460 14872 477466 14884
rect 488626 14872 488632 14884
rect 477460 14844 488632 14872
rect 477460 14832 477466 14844
rect 488626 14832 488632 14844
rect 488684 14832 488690 14884
rect 81434 14764 81440 14816
rect 81492 14804 81498 14816
rect 216858 14804 216864 14816
rect 81492 14776 216864 14804
rect 81492 14764 81498 14776
rect 216858 14764 216864 14776
rect 216916 14764 216922 14816
rect 233510 14764 233516 14816
rect 233568 14804 233574 14816
rect 242894 14804 242900 14816
rect 233568 14776 242900 14804
rect 233568 14764 233574 14776
rect 242894 14764 242900 14776
rect 242952 14764 242958 14816
rect 244550 14764 244556 14816
rect 244608 14804 244614 14816
rect 284478 14804 284484 14816
rect 244608 14776 284484 14804
rect 244608 14764 244614 14776
rect 284478 14764 284484 14776
rect 284536 14764 284542 14816
rect 295334 14764 295340 14816
rect 295392 14804 295398 14816
rect 407114 14804 407120 14816
rect 295392 14776 407120 14804
rect 295392 14764 295398 14776
rect 407114 14764 407120 14776
rect 407172 14764 407178 14816
rect 412634 14764 412640 14816
rect 412692 14804 412698 14816
rect 423582 14804 423588 14816
rect 412692 14776 423588 14804
rect 412692 14764 412698 14776
rect 423582 14764 423588 14776
rect 423640 14764 423646 14816
rect 423674 14764 423680 14816
rect 423732 14804 423738 14816
rect 435818 14804 435824 14816
rect 423732 14776 435824 14804
rect 423732 14764 423738 14776
rect 435818 14764 435824 14776
rect 435876 14764 435882 14816
rect 439222 14764 439228 14816
rect 439280 14804 439286 14816
rect 445110 14804 445116 14816
rect 439280 14776 445116 14804
rect 439280 14764 439286 14776
rect 445110 14764 445116 14776
rect 445168 14764 445174 14816
rect 448698 14764 448704 14816
rect 448756 14804 448762 14816
rect 513282 14804 513288 14816
rect 448756 14776 513288 14804
rect 448756 14764 448762 14776
rect 513282 14764 513288 14776
rect 513340 14764 513346 14816
rect 69842 14696 69848 14748
rect 69900 14736 69906 14748
rect 78306 14736 78312 14748
rect 69900 14708 78312 14736
rect 69900 14696 69906 14708
rect 78306 14696 78312 14708
rect 78364 14696 78370 14748
rect 81894 14696 81900 14748
rect 81952 14736 81958 14748
rect 223022 14736 223028 14748
rect 81952 14708 223028 14736
rect 81952 14696 81958 14708
rect 223022 14696 223028 14708
rect 223080 14696 223086 14748
rect 223482 14696 223488 14748
rect 223540 14736 223546 14748
rect 317966 14736 317972 14748
rect 223540 14708 317972 14736
rect 223540 14696 223546 14708
rect 317966 14696 317972 14708
rect 318024 14696 318030 14748
rect 322750 14696 322756 14748
rect 322808 14736 322814 14748
rect 450906 14736 450912 14748
rect 322808 14708 450912 14736
rect 322808 14696 322814 14708
rect 450906 14696 450912 14708
rect 450964 14696 450970 14748
rect 460290 14696 460296 14748
rect 460348 14736 460354 14748
rect 471238 14736 471244 14748
rect 460348 14708 471244 14736
rect 460348 14696 460354 14708
rect 471238 14696 471244 14708
rect 471296 14696 471302 14748
rect 480254 14696 480260 14748
rect 480312 14736 480318 14748
rect 507210 14736 507216 14748
rect 480312 14708 507216 14736
rect 480312 14696 480318 14708
rect 507210 14696 507216 14708
rect 507268 14696 507274 14748
rect 65582 14640 70394 14668
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 21450 14600 21456 14612
rect 5316 14572 21456 14600
rect 5316 14560 5322 14572
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 22370 14560 22376 14612
rect 22428 14600 22434 14612
rect 47302 14600 47308 14612
rect 22428 14572 47308 14600
rect 22428 14560 22434 14572
rect 47302 14560 47308 14572
rect 47360 14560 47366 14612
rect 57054 14560 57060 14612
rect 57112 14600 57118 14612
rect 60090 14600 60096 14612
rect 57112 14572 60096 14600
rect 57112 14560 57118 14572
rect 60090 14560 60096 14572
rect 60148 14560 60154 14612
rect 64230 14560 64236 14612
rect 64288 14600 64294 14612
rect 67726 14600 67732 14612
rect 64288 14572 67732 14600
rect 64288 14560 64294 14572
rect 67726 14560 67732 14572
rect 67784 14560 67790 14612
rect 70366 14600 70394 14640
rect 76374 14628 76380 14680
rect 76432 14668 76438 14680
rect 234614 14668 234620 14680
rect 76432 14640 234620 14668
rect 76432 14628 76438 14640
rect 234614 14628 234620 14640
rect 234672 14628 234678 14680
rect 240502 14628 240508 14680
rect 240560 14668 240566 14680
rect 396074 14668 396080 14680
rect 240560 14640 396080 14668
rect 240560 14628 240566 14640
rect 396074 14628 396080 14640
rect 396132 14628 396138 14680
rect 406562 14628 406568 14680
rect 406620 14668 406626 14680
rect 427078 14668 427084 14680
rect 406620 14640 427084 14668
rect 406620 14628 406626 14640
rect 427078 14628 427084 14640
rect 427136 14628 427142 14680
rect 427630 14628 427636 14680
rect 427688 14668 427694 14680
rect 493318 14668 493324 14680
rect 427688 14640 493324 14668
rect 427688 14628 427694 14640
rect 493318 14628 493324 14640
rect 493376 14628 493382 14680
rect 79134 14600 79140 14612
rect 70366 14572 79140 14600
rect 79134 14560 79140 14572
rect 79192 14560 79198 14612
rect 86126 14560 86132 14612
rect 86184 14600 86190 14612
rect 297266 14600 297272 14612
rect 86184 14572 297272 14600
rect 86184 14560 86190 14572
rect 297266 14560 297272 14572
rect 297324 14560 297330 14612
rect 355962 14560 355968 14612
rect 356020 14600 356026 14612
rect 521654 14600 521660 14612
rect 356020 14572 521660 14600
rect 356020 14560 356026 14572
rect 521654 14560 521660 14572
rect 521712 14560 521718 14612
rect 1026 14492 1032 14544
rect 1084 14532 1090 14544
rect 13814 14532 13820 14544
rect 1084 14504 13820 14532
rect 1084 14492 1090 14504
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 17034 14492 17040 14544
rect 17092 14532 17098 14544
rect 42518 14532 42524 14544
rect 17092 14504 42524 14532
rect 17092 14492 17098 14504
rect 42518 14492 42524 14504
rect 42576 14492 42582 14544
rect 54110 14492 54116 14544
rect 54168 14532 54174 14544
rect 79226 14532 79232 14544
rect 54168 14504 79232 14532
rect 54168 14492 54174 14504
rect 79226 14492 79232 14504
rect 79284 14492 79290 14544
rect 89070 14492 89076 14544
rect 89128 14532 89134 14544
rect 282178 14532 282184 14544
rect 89128 14504 282184 14532
rect 89128 14492 89134 14504
rect 282178 14492 282184 14504
rect 282236 14492 282242 14544
rect 283374 14492 283380 14544
rect 283432 14532 283438 14544
rect 498930 14532 498936 14544
rect 283432 14504 498936 14532
rect 283432 14492 283438 14504
rect 498930 14492 498936 14504
rect 498988 14492 498994 14544
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 40218 14464 40224 14476
rect 2924 14436 40224 14464
rect 2924 14424 2930 14436
rect 40218 14424 40224 14436
rect 40276 14424 40282 14476
rect 40310 14424 40316 14476
rect 40368 14464 40374 14476
rect 40678 14464 40684 14476
rect 40368 14436 40684 14464
rect 40368 14424 40374 14436
rect 40678 14424 40684 14436
rect 40736 14424 40742 14476
rect 55214 14424 55220 14476
rect 55272 14464 55278 14476
rect 79502 14464 79508 14476
rect 55272 14436 79508 14464
rect 55272 14424 55278 14436
rect 79502 14424 79508 14436
rect 79560 14424 79566 14476
rect 81526 14424 81532 14476
rect 81584 14464 81590 14476
rect 251818 14464 251824 14476
rect 81584 14436 251824 14464
rect 81584 14424 81590 14436
rect 251818 14424 251824 14436
rect 251876 14424 251882 14476
rect 263134 14424 263140 14476
rect 263192 14464 263198 14476
rect 570322 14464 570328 14476
rect 263192 14436 570328 14464
rect 263192 14424 263198 14436
rect 570322 14424 570328 14436
rect 570380 14424 570386 14476
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 21082 14396 21088 14408
rect 9180 14368 21088 14396
rect 9180 14356 9186 14368
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 30834 14356 30840 14408
rect 30892 14396 30898 14408
rect 44726 14396 44732 14408
rect 30892 14368 44732 14396
rect 30892 14356 30898 14368
rect 44726 14356 44732 14368
rect 44784 14356 44790 14408
rect 60366 14356 60372 14408
rect 60424 14396 60430 14408
rect 131298 14396 131304 14408
rect 60424 14368 131304 14396
rect 60424 14356 60430 14368
rect 131298 14356 131304 14368
rect 131356 14356 131362 14408
rect 445018 14356 445024 14408
rect 445076 14396 445082 14408
rect 448514 14396 448520 14408
rect 445076 14368 448520 14396
rect 445076 14356 445082 14368
rect 448514 14356 448520 14368
rect 448572 14356 448578 14408
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 21266 14328 21272 14340
rect 15712 14300 21272 14328
rect 15712 14288 15718 14300
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 61286 14288 61292 14340
rect 61344 14328 61350 14340
rect 108298 14328 108304 14340
rect 61344 14300 108304 14328
rect 61344 14288 61350 14300
rect 108298 14288 108304 14300
rect 108356 14288 108362 14340
rect 64690 14220 64696 14272
rect 64748 14260 64754 14272
rect 88242 14260 88248 14272
rect 64748 14232 88248 14260
rect 64748 14220 64754 14232
rect 88242 14220 88248 14232
rect 88300 14220 88306 14272
rect 93578 14220 93584 14272
rect 93636 14260 93642 14272
rect 97534 14260 97540 14272
rect 93636 14232 97540 14260
rect 93636 14220 93642 14232
rect 97534 14220 97540 14232
rect 97592 14220 97598 14272
rect 441982 14220 441988 14272
rect 442040 14260 442046 14272
rect 448606 14260 448612 14272
rect 442040 14232 448612 14260
rect 442040 14220 442046 14232
rect 448606 14220 448612 14232
rect 448664 14220 448670 14272
rect 50798 14152 50804 14204
rect 50856 14192 50862 14204
rect 69842 14192 69848 14204
rect 50856 14164 69848 14192
rect 50856 14152 50862 14164
rect 69842 14152 69848 14164
rect 69900 14152 69906 14204
rect 79226 14152 79232 14204
rect 79284 14192 79290 14204
rect 84930 14192 84936 14204
rect 79284 14164 84936 14192
rect 79284 14152 79290 14164
rect 84930 14152 84936 14164
rect 84988 14152 84994 14204
rect 168558 14192 168564 14204
rect 85592 14164 168564 14192
rect 58710 14084 58716 14136
rect 58768 14124 58774 14136
rect 77202 14124 77208 14136
rect 58768 14096 77208 14124
rect 58768 14084 58774 14096
rect 77202 14084 77208 14096
rect 77260 14084 77266 14136
rect 79686 14084 79692 14136
rect 79744 14124 79750 14136
rect 85592 14124 85620 14164
rect 168558 14152 168564 14164
rect 168616 14152 168622 14204
rect 420914 14152 420920 14204
rect 420972 14192 420978 14204
rect 424962 14192 424968 14204
rect 420972 14164 424968 14192
rect 420972 14152 420978 14164
rect 424962 14152 424968 14164
rect 425020 14152 425026 14204
rect 79744 14096 85620 14124
rect 79744 14084 79750 14096
rect 93486 14084 93492 14136
rect 93544 14124 93550 14136
rect 148962 14124 148968 14136
rect 93544 14096 148968 14124
rect 93544 14084 93550 14096
rect 148962 14084 148968 14096
rect 149020 14084 149026 14136
rect 417418 14084 417424 14136
rect 417476 14124 417482 14136
rect 423766 14124 423772 14136
rect 417476 14096 423772 14124
rect 417476 14084 417482 14096
rect 423766 14084 423772 14096
rect 423824 14084 423830 14136
rect 66530 14016 66536 14068
rect 66588 14056 66594 14068
rect 81434 14056 81440 14068
rect 66588 14028 81440 14056
rect 66588 14016 66594 14028
rect 81434 14016 81440 14028
rect 81492 14016 81498 14068
rect 108482 14016 108488 14068
rect 108540 14056 108546 14068
rect 113634 14056 113640 14068
rect 108540 14028 113640 14056
rect 108540 14016 108546 14028
rect 113634 14016 113640 14028
rect 113692 14016 113698 14068
rect 117682 14016 117688 14068
rect 117740 14056 117746 14068
rect 119890 14056 119896 14068
rect 117740 14028 119896 14056
rect 117740 14016 117746 14028
rect 119890 14016 119896 14028
rect 119948 14016 119954 14068
rect 157334 14016 157340 14068
rect 157392 14056 157398 14068
rect 159542 14056 159548 14068
rect 157392 14028 159548 14056
rect 157392 14016 157398 14028
rect 159542 14016 159548 14028
rect 159600 14016 159606 14068
rect 78950 13948 78956 14000
rect 79008 13988 79014 14000
rect 80882 13988 80888 14000
rect 79008 13960 80888 13988
rect 79008 13948 79014 13960
rect 80882 13948 80888 13960
rect 80940 13948 80946 14000
rect 82170 13948 82176 14000
rect 82228 13988 82234 14000
rect 188522 13988 188528 14000
rect 82228 13960 188528 13988
rect 82228 13948 82234 13960
rect 188522 13948 188528 13960
rect 188580 13948 188586 14000
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 92382 13920 92388 13932
rect 19024 13892 92388 13920
rect 19024 13880 19030 13892
rect 92382 13880 92388 13892
rect 92440 13880 92446 13932
rect 115934 13880 115940 13932
rect 115992 13920 115998 13932
rect 117958 13920 117964 13932
rect 115992 13892 117964 13920
rect 115992 13880 115998 13892
rect 117958 13880 117964 13892
rect 118016 13880 118022 13932
rect 118786 13880 118792 13932
rect 118844 13920 118850 13932
rect 121730 13920 121736 13932
rect 118844 13892 121736 13920
rect 118844 13880 118850 13892
rect 121730 13880 121736 13892
rect 121788 13880 121794 13932
rect 123294 13880 123300 13932
rect 123352 13920 123358 13932
rect 129734 13920 129740 13932
rect 123352 13892 129740 13920
rect 123352 13880 123358 13892
rect 129734 13880 129740 13892
rect 129792 13880 129798 13932
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 19334 13852 19340 13864
rect 18196 13824 19340 13852
rect 18196 13812 18202 13824
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 27614 13812 27620 13864
rect 27672 13852 27678 13864
rect 33870 13852 33876 13864
rect 27672 13824 33876 13852
rect 27672 13812 27678 13824
rect 33870 13812 33876 13824
rect 33928 13812 33934 13864
rect 78674 13812 78680 13864
rect 78732 13852 78738 13864
rect 81986 13852 81992 13864
rect 78732 13824 81992 13852
rect 78732 13812 78738 13824
rect 81986 13812 81992 13824
rect 82044 13812 82050 13864
rect 102134 13812 102140 13864
rect 102192 13852 102198 13864
rect 108114 13852 108120 13864
rect 102192 13824 108120 13852
rect 102192 13812 102198 13824
rect 108114 13812 108120 13824
rect 108172 13812 108178 13864
rect 108298 13812 108304 13864
rect 108356 13852 108362 13864
rect 125502 13852 125508 13864
rect 108356 13824 125508 13852
rect 108356 13812 108362 13824
rect 125502 13812 125508 13824
rect 125560 13812 125566 13864
rect 126514 13812 126520 13864
rect 126572 13852 126578 13864
rect 127618 13852 127624 13864
rect 126572 13824 127624 13852
rect 126572 13812 126578 13824
rect 127618 13812 127624 13824
rect 127676 13812 127682 13864
rect 137278 13852 137284 13864
rect 132466 13824 137284 13852
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 10962 13784 10968 13796
rect 5408 13756 10968 13784
rect 5408 13744 5414 13756
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 65702 13784 65708 13796
rect 12406 13756 65708 13784
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 12406 13716 12434 13756
rect 65702 13744 65708 13756
rect 65760 13744 65766 13796
rect 67634 13744 67640 13796
rect 67692 13784 67698 13796
rect 71774 13784 71780 13796
rect 67692 13756 71780 13784
rect 67692 13744 67698 13756
rect 71774 13744 71780 13756
rect 71832 13744 71838 13796
rect 83182 13744 83188 13796
rect 83240 13784 83246 13796
rect 86770 13784 86776 13796
rect 83240 13756 86776 13784
rect 83240 13744 83246 13756
rect 86770 13744 86776 13756
rect 86828 13744 86834 13796
rect 114554 13744 114560 13796
rect 114612 13784 114618 13796
rect 118786 13784 118792 13796
rect 114612 13756 118792 13784
rect 114612 13744 114618 13756
rect 118786 13744 118792 13756
rect 118844 13744 118850 13796
rect 122190 13744 122196 13796
rect 122248 13784 122254 13796
rect 132466 13784 132494 13824
rect 137278 13812 137284 13824
rect 137336 13812 137342 13864
rect 149054 13812 149060 13864
rect 149112 13852 149118 13864
rect 152734 13852 152740 13864
rect 149112 13824 152740 13852
rect 149112 13812 149118 13824
rect 152734 13812 152740 13824
rect 152792 13812 152798 13864
rect 435542 13812 435548 13864
rect 435600 13852 435606 13864
rect 440878 13852 440884 13864
rect 435600 13824 440884 13852
rect 435600 13812 435606 13824
rect 440878 13812 440884 13824
rect 440936 13812 440942 13864
rect 122248 13756 132494 13784
rect 122248 13744 122254 13756
rect 155954 13744 155960 13796
rect 156012 13784 156018 13796
rect 159450 13784 159456 13796
rect 156012 13756 159456 13784
rect 156012 13744 156018 13756
rect 159450 13744 159456 13756
rect 159508 13744 159514 13796
rect 201402 13744 201408 13796
rect 201460 13784 201466 13796
rect 327534 13784 327540 13796
rect 201460 13756 327540 13784
rect 201460 13744 201466 13756
rect 327534 13744 327540 13756
rect 327592 13744 327598 13796
rect 4028 13688 12434 13716
rect 4028 13676 4034 13688
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 66438 13716 66444 13728
rect 13872 13688 66444 13716
rect 13872 13676 13878 13688
rect 66438 13676 66444 13688
rect 66496 13676 66502 13728
rect 75270 13676 75276 13728
rect 75328 13716 75334 13728
rect 211798 13716 211804 13728
rect 75328 13688 211804 13716
rect 75328 13676 75334 13688
rect 211798 13676 211804 13688
rect 211856 13676 211862 13728
rect 15470 13608 15476 13660
rect 15528 13648 15534 13660
rect 67818 13648 67824 13660
rect 15528 13620 67824 13648
rect 15528 13608 15534 13620
rect 67818 13608 67824 13620
rect 67876 13608 67882 13660
rect 73062 13608 73068 13660
rect 73120 13648 73126 13660
rect 211062 13648 211068 13660
rect 73120 13620 211068 13648
rect 73120 13608 73126 13620
rect 211062 13608 211068 13620
rect 211120 13608 211126 13660
rect 223022 13608 223028 13660
rect 223080 13648 223086 13660
rect 241422 13648 241428 13660
rect 223080 13620 241428 13648
rect 223080 13608 223086 13620
rect 241422 13608 241428 13620
rect 241480 13608 241486 13660
rect 18230 13540 18236 13592
rect 18288 13580 18294 13592
rect 68370 13580 68376 13592
rect 18288 13552 68376 13580
rect 18288 13540 18294 13552
rect 68370 13540 68376 13552
rect 68428 13540 68434 13592
rect 78490 13540 78496 13592
rect 78548 13580 78554 13592
rect 229370 13580 229376 13592
rect 78548 13552 229376 13580
rect 78548 13540 78554 13552
rect 229370 13540 229376 13552
rect 229428 13540 229434 13592
rect 10318 13472 10324 13524
rect 10376 13512 10382 13524
rect 23658 13512 23664 13524
rect 10376 13484 23664 13512
rect 10376 13472 10382 13484
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 33502 13472 33508 13524
rect 33560 13512 33566 13524
rect 37182 13512 37188 13524
rect 33560 13484 37188 13512
rect 33560 13472 33566 13484
rect 37182 13472 37188 13484
rect 37240 13472 37246 13524
rect 53742 13472 53748 13524
rect 53800 13512 53806 13524
rect 57330 13512 57336 13524
rect 53800 13484 57336 13512
rect 53800 13472 53806 13484
rect 57330 13472 57336 13484
rect 57388 13472 57394 13524
rect 81158 13472 81164 13524
rect 81216 13512 81222 13524
rect 255314 13512 255320 13524
rect 81216 13484 255320 13512
rect 81216 13472 81222 13484
rect 255314 13472 255320 13484
rect 255372 13472 255378 13524
rect 276014 13472 276020 13524
rect 276072 13512 276078 13524
rect 282914 13512 282920 13524
rect 276072 13484 282920 13512
rect 276072 13472 276078 13484
rect 282914 13472 282920 13484
rect 282972 13472 282978 13524
rect 31662 13404 31668 13456
rect 31720 13444 31726 13456
rect 36814 13444 36820 13456
rect 31720 13416 36820 13444
rect 31720 13404 31726 13416
rect 36814 13404 36820 13416
rect 36872 13404 36878 13456
rect 65794 13404 65800 13456
rect 65852 13444 65858 13456
rect 70394 13444 70400 13456
rect 65852 13416 70400 13444
rect 65852 13404 65858 13416
rect 70394 13404 70400 13416
rect 70452 13404 70458 13456
rect 89898 13404 89904 13456
rect 89956 13444 89962 13456
rect 244274 13444 244280 13456
rect 89956 13416 244280 13444
rect 89956 13404 89962 13416
rect 244274 13404 244280 13416
rect 244332 13404 244338 13456
rect 253934 13404 253940 13456
rect 253992 13444 253998 13456
rect 432046 13444 432052 13456
rect 253992 13416 432052 13444
rect 253992 13404 253998 13416
rect 432046 13404 432052 13416
rect 432104 13404 432110 13456
rect 21818 13336 21824 13388
rect 21876 13376 21882 13388
rect 43254 13376 43260 13388
rect 21876 13348 43260 13376
rect 21876 13336 21882 13348
rect 43254 13336 43260 13348
rect 43312 13336 43318 13388
rect 50982 13336 50988 13388
rect 51040 13376 51046 13388
rect 70946 13376 70952 13388
rect 51040 13348 70952 13376
rect 51040 13336 51046 13348
rect 70946 13336 70952 13348
rect 71004 13336 71010 13388
rect 80790 13336 80796 13388
rect 80848 13376 80854 13388
rect 258718 13376 258724 13388
rect 80848 13348 258724 13376
rect 80848 13336 80854 13348
rect 258718 13336 258724 13348
rect 258776 13336 258782 13388
rect 282178 13336 282184 13388
rect 282236 13376 282242 13388
rect 314010 13376 314016 13388
rect 282236 13348 314016 13376
rect 282236 13336 282242 13348
rect 314010 13336 314016 13348
rect 314068 13336 314074 13388
rect 363598 13336 363604 13388
rect 363656 13376 363662 13388
rect 398926 13376 398932 13388
rect 363656 13348 398932 13376
rect 363656 13336 363662 13348
rect 398926 13336 398932 13348
rect 398984 13336 398990 13388
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 40034 13308 40040 13320
rect 18012 13280 40040 13308
rect 18012 13268 18018 13280
rect 40034 13268 40040 13280
rect 40092 13268 40098 13320
rect 51534 13268 51540 13320
rect 51592 13308 51598 13320
rect 74994 13308 75000 13320
rect 51592 13280 75000 13308
rect 51592 13268 51598 13280
rect 74994 13268 75000 13280
rect 75052 13268 75058 13320
rect 86678 13268 86684 13320
rect 86736 13308 86742 13320
rect 276014 13308 276020 13320
rect 86736 13280 276020 13308
rect 86736 13268 86742 13280
rect 276014 13268 276020 13280
rect 276072 13268 276078 13320
rect 280338 13268 280344 13320
rect 280396 13308 280402 13320
rect 285766 13308 285772 13320
rect 280396 13280 285772 13308
rect 280396 13268 280402 13280
rect 285766 13268 285772 13280
rect 285824 13268 285830 13320
rect 298462 13268 298468 13320
rect 298520 13308 298526 13320
rect 405826 13308 405832 13320
rect 298520 13280 405832 13308
rect 298520 13268 298526 13280
rect 405826 13268 405832 13280
rect 405884 13268 405890 13320
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 40586 13240 40592 13252
rect 13688 13212 40592 13240
rect 13688 13200 13694 13212
rect 40586 13200 40592 13212
rect 40644 13200 40650 13252
rect 54662 13200 54668 13252
rect 54720 13240 54726 13252
rect 82170 13240 82176 13252
rect 54720 13212 82176 13240
rect 54720 13200 54726 13212
rect 82170 13200 82176 13212
rect 82228 13200 82234 13252
rect 91554 13200 91560 13252
rect 91612 13240 91618 13252
rect 307846 13240 307852 13252
rect 91612 13212 307852 13240
rect 91612 13200 91618 13212
rect 307846 13200 307852 13212
rect 307904 13200 307910 13252
rect 318058 13200 318064 13252
rect 318116 13240 318122 13252
rect 520274 13240 520280 13252
rect 318116 13212 520280 13240
rect 318116 13200 318122 13212
rect 520274 13200 520280 13212
rect 520332 13200 520338 13252
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 79226 13172 79232 13184
rect 17000 13144 79232 13172
rect 17000 13132 17006 13144
rect 79226 13132 79232 13144
rect 79284 13132 79290 13184
rect 91646 13132 91652 13184
rect 91704 13172 91710 13184
rect 318610 13172 318616 13184
rect 91704 13144 318616 13172
rect 91704 13132 91710 13144
rect 318610 13132 318616 13144
rect 318668 13132 318674 13184
rect 319530 13132 319536 13184
rect 319588 13172 319594 13184
rect 351914 13172 351920 13184
rect 319588 13144 351920 13172
rect 319588 13132 319594 13144
rect 351914 13132 351920 13144
rect 351972 13132 351978 13184
rect 355318 13132 355324 13184
rect 355376 13172 355382 13184
rect 417234 13172 417240 13184
rect 355376 13144 417240 13172
rect 355376 13132 355382 13144
rect 417234 13132 417240 13144
rect 417292 13132 417298 13184
rect 3878 13064 3884 13116
rect 3936 13104 3942 13116
rect 23474 13104 23480 13116
rect 3936 13076 23480 13104
rect 3936 13064 3942 13076
rect 23474 13064 23480 13076
rect 23532 13064 23538 13116
rect 24854 13064 24860 13116
rect 24912 13104 24918 13116
rect 33134 13104 33140 13116
rect 24912 13076 33140 13104
rect 24912 13064 24918 13076
rect 33134 13064 33140 13076
rect 33192 13064 33198 13116
rect 33686 13064 33692 13116
rect 33744 13104 33750 13116
rect 68830 13104 68836 13116
rect 33744 13076 68836 13104
rect 33744 13064 33750 13076
rect 68830 13064 68836 13076
rect 68888 13064 68894 13116
rect 77478 13064 77484 13116
rect 77536 13104 77542 13116
rect 241698 13104 241704 13116
rect 77536 13076 241704 13104
rect 77536 13064 77542 13076
rect 241698 13064 241704 13076
rect 241756 13064 241762 13116
rect 243538 13064 243544 13116
rect 243596 13104 243602 13116
rect 516134 13104 516140 13116
rect 243596 13076 516140 13104
rect 243596 13064 243602 13076
rect 516134 13064 516140 13076
rect 516192 13064 516198 13116
rect 11974 12996 11980 13048
rect 12032 13036 12038 13048
rect 21358 13036 21364 13048
rect 12032 13008 21364 13036
rect 12032 12996 12038 13008
rect 21358 12996 21364 13008
rect 21416 12996 21422 13048
rect 68738 12996 68744 13048
rect 68796 13036 68802 13048
rect 168374 13036 168380 13048
rect 68796 13008 168380 13036
rect 68796 12996 68802 13008
rect 168374 12996 168380 13008
rect 168432 12996 168438 13048
rect 210970 12996 210976 13048
rect 211028 13036 211034 13048
rect 299382 13036 299388 13048
rect 211028 13008 299388 13036
rect 211028 12996 211034 13008
rect 299382 12996 299388 13008
rect 299440 12996 299446 13048
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 91186 12968 91192 12980
rect 9364 12940 91192 12968
rect 9364 12928 9370 12940
rect 91186 12928 91192 12940
rect 91244 12928 91250 12980
rect 108114 12928 108120 12980
rect 108172 12968 108178 12980
rect 119430 12968 119436 12980
rect 108172 12940 119436 12968
rect 108172 12928 108178 12940
rect 119430 12928 119436 12940
rect 119488 12928 119494 12980
rect 119522 12928 119528 12980
rect 119580 12968 119586 12980
rect 156782 12968 156788 12980
rect 119580 12940 156788 12968
rect 119580 12928 119586 12940
rect 156782 12928 156788 12940
rect 156840 12928 156846 12980
rect 168558 12928 168564 12980
rect 168616 12968 168622 12980
rect 222102 12968 222108 12980
rect 168616 12940 222108 12968
rect 168616 12928 168622 12940
rect 222102 12928 222108 12940
rect 222160 12928 222166 12980
rect 58526 12860 58532 12912
rect 58584 12900 58590 12912
rect 115842 12900 115848 12912
rect 58584 12872 115848 12900
rect 58584 12860 58590 12872
rect 115842 12860 115848 12872
rect 115900 12860 115906 12912
rect 118050 12860 118056 12912
rect 118108 12900 118114 12912
rect 118418 12900 118424 12912
rect 118108 12872 118424 12900
rect 118108 12860 118114 12872
rect 118418 12860 118424 12872
rect 118476 12860 118482 12912
rect 84654 12792 84660 12844
rect 84712 12832 84718 12844
rect 87966 12832 87972 12844
rect 84712 12804 87972 12832
rect 84712 12792 84718 12804
rect 87966 12792 87972 12804
rect 88024 12792 88030 12844
rect 59078 12724 59084 12776
rect 59136 12764 59142 12776
rect 102134 12764 102140 12776
rect 59136 12736 102140 12764
rect 59136 12724 59142 12736
rect 102134 12724 102140 12736
rect 102192 12724 102198 12776
rect 70854 12656 70860 12708
rect 70912 12696 70918 12708
rect 179414 12696 179420 12708
rect 70912 12668 179420 12696
rect 70912 12656 70918 12668
rect 179414 12656 179420 12668
rect 179472 12656 179478 12708
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 91094 12628 91100 12640
rect 8260 12600 91100 12628
rect 8260 12588 8266 12600
rect 91094 12588 91100 12600
rect 91152 12588 91158 12640
rect 133782 12520 133788 12572
rect 133840 12560 133846 12572
rect 140130 12560 140136 12572
rect 133840 12532 140136 12560
rect 133840 12520 133846 12532
rect 140130 12520 140136 12532
rect 140188 12520 140194 12572
rect 89530 12452 89536 12504
rect 89588 12492 89594 12504
rect 90634 12492 90640 12504
rect 89588 12464 90640 12492
rect 89588 12452 89594 12464
rect 90634 12452 90640 12464
rect 90692 12452 90698 12504
rect 93688 12464 93992 12492
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 93688 12424 93716 12464
rect 8076 12396 93716 12424
rect 93964 12424 93992 12464
rect 102134 12452 102140 12504
rect 102192 12492 102198 12504
rect 105630 12492 105636 12504
rect 102192 12464 105636 12492
rect 102192 12452 102198 12464
rect 105630 12452 105636 12464
rect 105688 12452 105694 12504
rect 96430 12424 96436 12436
rect 93964 12396 96436 12424
rect 8076 12384 8082 12396
rect 96430 12384 96436 12396
rect 96488 12384 96494 12436
rect 106366 12384 106372 12436
rect 106424 12424 106430 12436
rect 116762 12424 116768 12436
rect 106424 12396 116768 12424
rect 106424 12384 106430 12396
rect 116762 12384 116768 12396
rect 116820 12384 116826 12436
rect 148318 12384 148324 12436
rect 148376 12424 148382 12436
rect 155862 12424 155868 12436
rect 148376 12396 155868 12424
rect 148376 12384 148382 12396
rect 155862 12384 155868 12396
rect 155920 12384 155926 12436
rect 168374 12384 168380 12436
rect 168432 12424 168438 12436
rect 180150 12424 180156 12436
rect 168432 12396 180156 12424
rect 168432 12384 168438 12396
rect 180150 12384 180156 12396
rect 180208 12384 180214 12436
rect 197354 12384 197360 12436
rect 197412 12424 197418 12436
rect 202690 12424 202696 12436
rect 197412 12396 202696 12424
rect 197412 12384 197418 12396
rect 202690 12384 202696 12396
rect 202748 12384 202754 12436
rect 377766 12384 377772 12436
rect 377824 12424 377830 12436
rect 380986 12424 380992 12436
rect 377824 12396 380992 12424
rect 377824 12384 377830 12396
rect 380986 12384 380992 12396
rect 381044 12384 381050 12436
rect 388530 12384 388536 12436
rect 388588 12424 388594 12436
rect 390922 12424 390928 12436
rect 388588 12396 390928 12424
rect 388588 12384 388594 12396
rect 390922 12384 390928 12396
rect 390980 12384 390986 12436
rect 403710 12384 403716 12436
rect 403768 12424 403774 12436
rect 408494 12424 408500 12436
rect 403768 12396 408500 12424
rect 403768 12384 403774 12396
rect 408494 12384 408500 12396
rect 408552 12384 408558 12436
rect 441614 12384 441620 12436
rect 441672 12424 441678 12436
rect 444650 12424 444656 12436
rect 441672 12396 444656 12424
rect 441672 12384 441678 12396
rect 444650 12384 444656 12396
rect 444708 12384 444714 12436
rect 1210 12316 1216 12368
rect 1268 12356 1274 12368
rect 69566 12356 69572 12368
rect 1268 12328 69572 12356
rect 1268 12316 1274 12328
rect 69566 12316 69572 12328
rect 69624 12316 69630 12368
rect 81434 12316 81440 12368
rect 81492 12356 81498 12368
rect 170306 12356 170312 12368
rect 81492 12328 170312 12356
rect 81492 12316 81498 12328
rect 170306 12316 170312 12328
rect 170364 12316 170370 12368
rect 423582 12316 423588 12368
rect 423640 12356 423646 12368
rect 435910 12356 435916 12368
rect 423640 12328 435916 12356
rect 423640 12316 423646 12328
rect 435910 12316 435916 12328
rect 435968 12316 435974 12368
rect 436002 12316 436008 12368
rect 436060 12356 436066 12368
rect 449802 12356 449808 12368
rect 436060 12328 449808 12356
rect 436060 12316 436066 12328
rect 449802 12316 449808 12328
rect 449860 12316 449866 12368
rect 2682 12248 2688 12300
rect 2740 12288 2746 12300
rect 67358 12288 67364 12300
rect 2740 12260 67364 12288
rect 2740 12248 2746 12260
rect 67358 12248 67364 12260
rect 67416 12248 67422 12300
rect 70302 12248 70308 12300
rect 70360 12288 70366 12300
rect 160186 12288 160192 12300
rect 70360 12260 160192 12288
rect 70360 12248 70366 12260
rect 160186 12248 160192 12260
rect 160244 12248 160250 12300
rect 179506 12248 179512 12300
rect 179564 12288 179570 12300
rect 241330 12288 241336 12300
rect 179564 12260 241336 12288
rect 179564 12248 179570 12260
rect 241330 12248 241336 12260
rect 241388 12248 241394 12300
rect 430574 12248 430580 12300
rect 430632 12288 430638 12300
rect 433978 12288 433984 12300
rect 430632 12260 433984 12288
rect 430632 12248 430638 12260
rect 433978 12248 433984 12260
rect 434036 12248 434042 12300
rect 442902 12248 442908 12300
rect 442960 12288 442966 12300
rect 448790 12288 448796 12300
rect 442960 12260 448796 12288
rect 442960 12248 442966 12260
rect 448790 12248 448796 12260
rect 448848 12248 448854 12300
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 24854 12220 24860 12232
rect 20588 12192 24860 12220
rect 20588 12180 20594 12192
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 72602 12180 72608 12232
rect 72660 12220 72666 12232
rect 183370 12220 183376 12232
rect 72660 12192 183376 12220
rect 72660 12180 72666 12192
rect 183370 12180 183376 12192
rect 183428 12180 183434 12232
rect 241422 12180 241428 12232
rect 241480 12220 241486 12232
rect 270034 12220 270040 12232
rect 241480 12192 270040 12220
rect 241480 12180 241486 12192
rect 270034 12180 270040 12192
rect 270092 12180 270098 12232
rect 417326 12180 417332 12232
rect 417384 12220 417390 12232
rect 443362 12220 443368 12232
rect 417384 12192 443368 12220
rect 417384 12180 417390 12192
rect 443362 12180 443368 12192
rect 443420 12180 443426 12232
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 12434 12152 12440 12164
rect 6880 12124 12440 12152
rect 6880 12112 6886 12124
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 21450 12112 21456 12164
rect 21508 12152 21514 12164
rect 23750 12152 23756 12164
rect 21508 12124 23756 12152
rect 21508 12112 21514 12124
rect 23750 12112 23756 12124
rect 23808 12112 23814 12164
rect 75822 12112 75828 12164
rect 75880 12152 75886 12164
rect 202230 12152 202236 12164
rect 75880 12124 202236 12152
rect 75880 12112 75886 12124
rect 202230 12112 202236 12124
rect 202288 12112 202294 12164
rect 222102 12112 222108 12164
rect 222160 12152 222166 12164
rect 255866 12152 255872 12164
rect 222160 12124 255872 12152
rect 222160 12112 222166 12124
rect 255866 12112 255872 12124
rect 255924 12112 255930 12164
rect 378042 12112 378048 12164
rect 378100 12152 378106 12164
rect 394970 12152 394976 12164
rect 378100 12124 394976 12152
rect 378100 12112 378106 12124
rect 394970 12112 394976 12124
rect 395028 12112 395034 12164
rect 427078 12112 427084 12164
rect 427136 12152 427142 12164
rect 463142 12152 463148 12164
rect 427136 12124 463148 12152
rect 427136 12112 427142 12124
rect 463142 12112 463148 12124
rect 463200 12112 463206 12164
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 19610 12084 19616 12096
rect 10652 12056 19616 12084
rect 10652 12044 10658 12056
rect 19610 12044 19616 12056
rect 19668 12044 19674 12096
rect 20898 12044 20904 12096
rect 20956 12084 20962 12096
rect 78674 12084 78680 12096
rect 20956 12056 78680 12084
rect 20956 12044 20962 12056
rect 78674 12044 78680 12056
rect 78732 12044 78738 12096
rect 85022 12044 85028 12096
rect 85080 12084 85086 12096
rect 223482 12084 223488 12096
rect 85080 12056 223488 12084
rect 85080 12044 85086 12056
rect 223482 12044 223488 12056
rect 223540 12044 223546 12096
rect 244274 12044 244280 12096
rect 244332 12084 244338 12096
rect 284570 12084 284576 12096
rect 244332 12056 284576 12084
rect 244332 12044 244338 12056
rect 284570 12044 284576 12056
rect 284628 12044 284634 12096
rect 395798 12044 395804 12096
rect 395856 12084 395862 12096
rect 395856 12056 441614 12084
rect 395856 12044 395862 12056
rect 10686 11976 10692 12028
rect 10744 12016 10750 12028
rect 20530 12016 20536 12028
rect 10744 11988 20536 12016
rect 10744 11976 10750 11988
rect 20530 11976 20536 11988
rect 20588 11976 20594 12028
rect 23474 11976 23480 12028
rect 23532 12016 23538 12028
rect 88794 12016 88800 12028
rect 23532 11988 88800 12016
rect 23532 11976 23538 11988
rect 88794 11976 88800 11988
rect 88852 11976 88858 12028
rect 88886 11976 88892 12028
rect 88944 12016 88950 12028
rect 93578 12016 93584 12028
rect 88944 11988 93584 12016
rect 88944 11976 88950 11988
rect 93578 11976 93584 11988
rect 93636 11976 93642 12028
rect 94682 11976 94688 12028
rect 94740 12016 94746 12028
rect 249702 12016 249708 12028
rect 94740 11988 249708 12016
rect 94740 11976 94746 11988
rect 249702 11976 249708 11988
rect 249760 11976 249766 12028
rect 255314 11976 255320 12028
rect 255372 12016 255378 12028
rect 264974 12016 264980 12028
rect 255372 11988 264980 12016
rect 255372 11976 255378 11988
rect 264974 11976 264980 11988
rect 265032 11976 265038 12028
rect 283006 11976 283012 12028
rect 283064 12016 283070 12028
rect 322198 12016 322204 12028
rect 283064 11988 322204 12016
rect 283064 11976 283070 11988
rect 322198 11976 322204 11988
rect 322256 11976 322262 12028
rect 358722 11976 358728 12028
rect 358780 12016 358786 12028
rect 434898 12016 434904 12028
rect 358780 11988 434904 12016
rect 358780 11976 358786 11988
rect 434898 11976 434904 11988
rect 434956 11976 434962 12028
rect 441586 12016 441614 12056
rect 448514 12044 448520 12096
rect 448572 12084 448578 12096
rect 460290 12084 460296 12096
rect 448572 12056 460296 12084
rect 448572 12044 448578 12056
rect 460290 12044 460296 12056
rect 460348 12044 460354 12096
rect 485038 12044 485044 12096
rect 485096 12084 485102 12096
rect 498286 12084 498292 12096
rect 485096 12056 498292 12084
rect 485096 12044 485102 12056
rect 498286 12044 498292 12056
rect 498344 12044 498350 12096
rect 448698 12016 448704 12028
rect 441586 11988 448704 12016
rect 448698 11976 448704 11988
rect 448756 11976 448762 12028
rect 448790 11976 448796 12028
rect 448848 12016 448854 12028
rect 459186 12016 459192 12028
rect 448848 11988 459192 12016
rect 448848 11976 448854 11988
rect 459186 11976 459192 11988
rect 459244 11976 459250 12028
rect 470594 11976 470600 12028
rect 470652 12016 470658 12028
rect 510246 12016 510252 12028
rect 470652 11988 510252 12016
rect 470652 11976 470658 11988
rect 510246 11976 510252 11988
rect 510304 11976 510310 12028
rect 8386 11908 8392 11960
rect 8444 11948 8450 11960
rect 18782 11948 18788 11960
rect 8444 11920 18788 11948
rect 8444 11908 8450 11920
rect 18782 11908 18788 11920
rect 18840 11908 18846 11960
rect 19058 11908 19064 11960
rect 19116 11948 19122 11960
rect 40678 11948 40684 11960
rect 19116 11920 40684 11948
rect 19116 11908 19122 11920
rect 40678 11908 40684 11920
rect 40736 11908 40742 11960
rect 55950 11908 55956 11960
rect 56008 11948 56014 11960
rect 66898 11948 66904 11960
rect 56008 11920 66904 11948
rect 56008 11908 56014 11920
rect 66898 11908 66904 11920
rect 66956 11908 66962 11960
rect 77202 11908 77208 11960
rect 77260 11948 77266 11960
rect 81526 11948 81532 11960
rect 77260 11920 81532 11948
rect 77260 11908 77266 11920
rect 81526 11908 81532 11920
rect 81584 11908 81590 11960
rect 82354 11908 82360 11960
rect 82412 11948 82418 11960
rect 245194 11948 245200 11960
rect 82412 11920 245200 11948
rect 82412 11908 82418 11920
rect 245194 11908 245200 11920
rect 245252 11908 245258 11960
rect 248506 11908 248512 11960
rect 248564 11948 248570 11960
rect 260650 11948 260656 11960
rect 248564 11920 260656 11948
rect 248564 11908 248570 11920
rect 260650 11908 260656 11920
rect 260708 11908 260714 11960
rect 262490 11908 262496 11960
rect 262548 11948 262554 11960
rect 348510 11948 348516 11960
rect 262548 11920 348516 11948
rect 262548 11908 262554 11920
rect 348510 11908 348516 11920
rect 348568 11908 348574 11960
rect 353294 11908 353300 11960
rect 353352 11948 353358 11960
rect 440234 11948 440240 11960
rect 353352 11920 440240 11948
rect 353352 11908 353358 11920
rect 440234 11908 440240 11920
rect 440292 11908 440298 11960
rect 448606 11908 448612 11960
rect 448664 11948 448670 11960
rect 491202 11948 491208 11960
rect 448664 11920 491208 11948
rect 448664 11908 448670 11920
rect 491202 11908 491208 11920
rect 491260 11908 491266 11960
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 41230 11880 41236 11892
rect 8812 11852 41236 11880
rect 8812 11840 8818 11852
rect 41230 11840 41236 11852
rect 41288 11840 41294 11892
rect 50430 11840 50436 11892
rect 50488 11880 50494 11892
rect 67634 11880 67640 11892
rect 50488 11852 67640 11880
rect 50488 11840 50494 11852
rect 67634 11840 67640 11852
rect 67692 11840 67698 11892
rect 82538 11840 82544 11892
rect 82596 11880 82602 11892
rect 261478 11880 261484 11892
rect 82596 11852 261484 11880
rect 82596 11840 82602 11852
rect 261478 11840 261484 11852
rect 261536 11840 261542 11892
rect 263594 11840 263600 11892
rect 263652 11880 263658 11892
rect 421558 11880 421564 11892
rect 263652 11852 421564 11880
rect 263652 11840 263658 11852
rect 421558 11840 421564 11852
rect 421616 11840 421622 11892
rect 435818 11840 435824 11892
rect 435876 11880 435882 11892
rect 488534 11880 488540 11892
rect 435876 11852 488540 11880
rect 435876 11840 435882 11852
rect 488534 11840 488540 11852
rect 488592 11840 488598 11892
rect 488626 11840 488632 11892
rect 488684 11880 488690 11892
rect 493962 11880 493968 11892
rect 488684 11852 493968 11880
rect 488684 11840 488690 11852
rect 493962 11840 493968 11852
rect 494020 11840 494026 11892
rect 63586 11812 63592 11824
rect 22940 11784 63592 11812
rect 1118 11704 1124 11756
rect 1176 11744 1182 11756
rect 15194 11744 15200 11756
rect 1176 11716 15200 11744
rect 1176 11704 1182 11716
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 18690 11704 18696 11756
rect 18748 11744 18754 11756
rect 22738 11744 22744 11756
rect 18748 11716 22744 11744
rect 18748 11704 18754 11716
rect 22738 11704 22744 11716
rect 22796 11704 22802 11756
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 22940 11676 22968 11784
rect 63586 11772 63592 11784
rect 63644 11772 63650 11824
rect 65518 11772 65524 11824
rect 65576 11812 65582 11824
rect 81342 11812 81348 11824
rect 65576 11784 81348 11812
rect 65576 11772 65582 11784
rect 81342 11772 81348 11784
rect 81400 11772 81406 11824
rect 88518 11772 88524 11824
rect 88576 11812 88582 11824
rect 303614 11812 303620 11824
rect 88576 11784 303620 11812
rect 88576 11772 88582 11784
rect 303614 11772 303620 11784
rect 303672 11772 303678 11824
rect 380894 11772 380900 11824
rect 380952 11812 380958 11824
rect 387794 11812 387800 11824
rect 380952 11784 387800 11812
rect 380952 11772 380958 11784
rect 387794 11772 387800 11784
rect 387852 11772 387858 11824
rect 390554 11772 390560 11824
rect 390612 11812 390618 11824
rect 520918 11812 520924 11824
rect 390612 11784 520924 11812
rect 390612 11772 390618 11784
rect 520918 11772 520924 11784
rect 520976 11772 520982 11824
rect 77202 11744 77208 11756
rect 18472 11648 22968 11676
rect 23032 11716 77208 11744
rect 18472 11636 18478 11648
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 22186 11608 22192 11620
rect 20220 11580 22192 11608
rect 20220 11568 20226 11580
rect 22186 11568 22192 11580
rect 22244 11568 22250 11620
rect 18874 11500 18880 11552
rect 18932 11540 18938 11552
rect 23032 11540 23060 11716
rect 77202 11704 77208 11716
rect 77260 11704 77266 11756
rect 79134 11704 79140 11756
rect 79192 11744 79198 11756
rect 93762 11744 93768 11756
rect 79192 11716 93768 11744
rect 79192 11704 79198 11716
rect 93762 11704 93768 11716
rect 93820 11704 93826 11756
rect 107838 11704 107844 11756
rect 107896 11744 107902 11756
rect 431402 11744 431408 11756
rect 107896 11716 431408 11744
rect 107896 11704 107902 11716
rect 431402 11704 431408 11716
rect 431460 11704 431466 11756
rect 438854 11704 438860 11756
rect 438912 11744 438918 11756
rect 445662 11744 445668 11756
rect 438912 11716 445668 11744
rect 438912 11704 438918 11716
rect 445662 11704 445668 11716
rect 445720 11704 445726 11756
rect 511994 11744 512000 11756
rect 451246 11716 512000 11744
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 43990 11676 43996 11688
rect 26292 11648 43996 11676
rect 26292 11636 26298 11648
rect 43990 11636 43996 11648
rect 44048 11636 44054 11688
rect 56870 11636 56876 11688
rect 56928 11676 56934 11688
rect 108390 11676 108396 11688
rect 56928 11648 108396 11676
rect 56928 11636 56934 11648
rect 108390 11636 108396 11648
rect 108448 11636 108454 11688
rect 218054 11636 218060 11688
rect 218112 11676 218118 11688
rect 219250 11676 219256 11688
rect 218112 11648 219256 11676
rect 218112 11636 218118 11648
rect 219250 11636 219256 11648
rect 219308 11636 219314 11688
rect 445478 11636 445484 11688
rect 445536 11676 445542 11688
rect 451246 11676 451274 11716
rect 511994 11704 512000 11716
rect 512052 11704 512058 11756
rect 513282 11704 513288 11756
rect 513340 11744 513346 11756
rect 531222 11744 531228 11756
rect 513340 11716 531228 11744
rect 513340 11704 513346 11716
rect 531222 11704 531228 11716
rect 531280 11704 531286 11756
rect 445536 11648 451274 11676
rect 445536 11636 445542 11648
rect 453298 11636 453304 11688
rect 453356 11676 453362 11688
rect 457438 11676 457444 11688
rect 453356 11648 457444 11676
rect 453356 11636 453362 11648
rect 457438 11636 457444 11648
rect 457496 11636 457502 11688
rect 480898 11636 480904 11688
rect 480956 11676 480962 11688
rect 485222 11676 485228 11688
rect 480956 11648 485228 11676
rect 480956 11636 480962 11648
rect 485222 11636 485228 11648
rect 485280 11636 485286 11688
rect 57790 11568 57796 11620
rect 57848 11608 57854 11620
rect 107010 11608 107016 11620
rect 57848 11580 107016 11608
rect 57848 11568 57854 11580
rect 107010 11568 107016 11580
rect 107068 11568 107074 11620
rect 18932 11512 23060 11540
rect 18932 11500 18938 11512
rect 58342 11500 58348 11552
rect 58400 11540 58406 11552
rect 82722 11540 82728 11552
rect 58400 11512 82728 11540
rect 58400 11500 58406 11512
rect 82722 11500 82728 11512
rect 82780 11500 82786 11552
rect 103698 11500 103704 11552
rect 103756 11540 103762 11552
rect 125134 11540 125140 11552
rect 103756 11512 125140 11540
rect 103756 11500 103762 11512
rect 125134 11500 125140 11512
rect 125192 11500 125198 11552
rect 15286 11432 15292 11484
rect 15344 11472 15350 11484
rect 71682 11472 71688 11484
rect 15344 11444 71688 11472
rect 15344 11432 15350 11444
rect 71682 11432 71688 11444
rect 71740 11432 71746 11484
rect 71774 11432 71780 11484
rect 71832 11472 71838 11484
rect 84562 11472 84568 11484
rect 71832 11444 84568 11472
rect 71832 11432 71838 11444
rect 84562 11432 84568 11444
rect 84620 11432 84626 11484
rect 95050 11432 95056 11484
rect 95108 11472 95114 11484
rect 110414 11472 110420 11484
rect 95108 11444 110420 11472
rect 95108 11432 95114 11444
rect 110414 11432 110420 11444
rect 110472 11432 110478 11484
rect 211062 11432 211068 11484
rect 211120 11472 211126 11484
rect 213362 11472 213368 11484
rect 211120 11444 213368 11472
rect 211120 11432 211126 11444
rect 213362 11432 213368 11444
rect 213420 11432 213426 11484
rect 67542 11364 67548 11416
rect 67600 11404 67606 11416
rect 151354 11404 151360 11416
rect 67600 11376 151360 11404
rect 67600 11364 67606 11376
rect 151354 11364 151360 11376
rect 151412 11364 151418 11416
rect 21266 11296 21272 11348
rect 21324 11336 21330 11348
rect 77018 11336 77024 11348
rect 21324 11308 77024 11336
rect 21324 11296 21330 11308
rect 77018 11296 77024 11308
rect 77076 11296 77082 11348
rect 133230 11296 133236 11348
rect 133288 11336 133294 11348
rect 136082 11336 136088 11348
rect 133288 11308 136088 11336
rect 133288 11296 133294 11308
rect 136082 11296 136088 11308
rect 136140 11296 136146 11348
rect 111794 11160 111800 11212
rect 111852 11200 111858 11212
rect 378042 11200 378048 11212
rect 111852 11172 378048 11200
rect 111852 11160 111858 11172
rect 378042 11160 378048 11172
rect 378100 11160 378106 11212
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 13504 11104 19288 11132
rect 13504 11092 13510 11104
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 10928 11036 19196 11064
rect 10928 11024 10934 11036
rect 19168 10928 19196 11036
rect 19260 10996 19288 11104
rect 116762 11092 116768 11144
rect 116820 11132 116826 11144
rect 398834 11132 398840 11144
rect 116820 11104 398840 11132
rect 116820 11092 116826 11104
rect 398834 11092 398840 11104
rect 398892 11092 398898 11144
rect 92934 11024 92940 11076
rect 92992 11064 92998 11076
rect 95050 11064 95056 11076
rect 92992 11036 95056 11064
rect 92992 11024 92998 11036
rect 95050 11024 95056 11036
rect 95108 11024 95114 11076
rect 95418 11024 95424 11076
rect 95476 11064 95482 11076
rect 97534 11064 97540 11076
rect 95476 11036 97540 11064
rect 95476 11024 95482 11036
rect 97534 11024 97540 11036
rect 97592 11024 97598 11076
rect 70578 10996 70584 11008
rect 19260 10968 70584 10996
rect 70578 10956 70584 10968
rect 70636 10956 70642 11008
rect 96890 10956 96896 11008
rect 96948 10996 96954 11008
rect 100754 10996 100760 11008
rect 96948 10968 100760 10996
rect 96948 10956 96954 10968
rect 100754 10956 100760 10968
rect 100812 10956 100818 11008
rect 106274 10956 106280 11008
rect 106332 10996 106338 11008
rect 107930 10996 107936 11008
rect 106332 10968 107936 10996
rect 106332 10956 106338 10968
rect 107930 10956 107936 10968
rect 107988 10956 107994 11008
rect 114094 10956 114100 11008
rect 114152 10996 114158 11008
rect 115842 10996 115848 11008
rect 114152 10968 115848 10996
rect 114152 10956 114158 10968
rect 115842 10956 115848 10968
rect 115900 10956 115906 11008
rect 151354 10956 151360 11008
rect 151412 10996 151418 11008
rect 151814 10996 151820 11008
rect 151412 10968 151820 10996
rect 151412 10956 151418 10968
rect 151814 10956 151820 10968
rect 151872 10956 151878 11008
rect 179414 10956 179420 11008
rect 179472 10996 179478 11008
rect 198734 10996 198740 11008
rect 179472 10968 198740 10996
rect 179472 10956 179478 10968
rect 198734 10956 198740 10968
rect 198792 10956 198798 11008
rect 19168 10900 20024 10928
rect 19996 10792 20024 10900
rect 59814 10888 59820 10940
rect 59872 10928 59878 10940
rect 61654 10928 61660 10940
rect 59872 10900 61660 10928
rect 59872 10888 59878 10900
rect 61654 10888 61660 10900
rect 61712 10888 61718 10940
rect 66162 10888 66168 10940
rect 66220 10928 66226 10940
rect 71130 10928 71136 10940
rect 66220 10900 71136 10928
rect 66220 10888 66226 10900
rect 71130 10888 71136 10900
rect 71188 10888 71194 10940
rect 78398 10888 78404 10940
rect 78456 10928 78462 10940
rect 183462 10928 183468 10940
rect 78456 10900 183468 10928
rect 78456 10888 78462 10900
rect 183462 10888 183468 10900
rect 183520 10888 183526 10940
rect 209866 10928 209872 10940
rect 190426 10900 209872 10928
rect 24854 10820 24860 10872
rect 24912 10860 24918 10872
rect 63126 10860 63132 10872
rect 24912 10832 63132 10860
rect 24912 10820 24918 10832
rect 63126 10820 63132 10832
rect 63184 10820 63190 10872
rect 68462 10820 68468 10872
rect 68520 10860 68526 10872
rect 182266 10860 182272 10872
rect 68520 10832 182272 10860
rect 68520 10820 68526 10832
rect 182266 10820 182272 10832
rect 182324 10820 182330 10872
rect 183370 10820 183376 10872
rect 183428 10860 183434 10872
rect 190426 10860 190454 10900
rect 209866 10888 209872 10900
rect 209924 10888 209930 10940
rect 210050 10888 210056 10940
rect 210108 10928 210114 10940
rect 235994 10928 236000 10940
rect 210108 10900 236000 10928
rect 210108 10888 210114 10900
rect 235994 10888 236000 10900
rect 236052 10888 236058 10940
rect 241330 10888 241336 10940
rect 241388 10928 241394 10940
rect 268378 10928 268384 10940
rect 241388 10900 268384 10928
rect 241388 10888 241394 10900
rect 268378 10888 268384 10900
rect 268436 10888 268442 10940
rect 276658 10928 276664 10940
rect 270696 10900 276664 10928
rect 183428 10832 190454 10860
rect 183428 10820 183434 10832
rect 223482 10820 223488 10872
rect 223540 10860 223546 10872
rect 270696 10860 270724 10900
rect 276658 10888 276664 10900
rect 276716 10888 276722 10940
rect 223540 10832 270724 10860
rect 223540 10820 223546 10832
rect 276014 10820 276020 10872
rect 276072 10860 276078 10872
rect 299474 10860 299480 10872
rect 276072 10832 299480 10860
rect 276072 10820 276078 10832
rect 299474 10820 299480 10832
rect 299532 10820 299538 10872
rect 85758 10792 85764 10804
rect 19996 10764 85764 10792
rect 85758 10752 85764 10764
rect 85816 10752 85822 10804
rect 88978 10752 88984 10804
rect 89036 10792 89042 10804
rect 223390 10792 223396 10804
rect 89036 10764 223396 10792
rect 89036 10752 89042 10764
rect 223390 10752 223396 10764
rect 223448 10752 223454 10804
rect 249702 10752 249708 10804
rect 249760 10792 249766 10804
rect 284294 10792 284300 10804
rect 249760 10764 284300 10792
rect 249760 10752 249766 10764
rect 284294 10752 284300 10764
rect 284352 10752 284358 10804
rect 303614 10752 303620 10804
rect 303672 10792 303678 10804
rect 312170 10792 312176 10804
rect 303672 10764 312176 10792
rect 303672 10752 303678 10764
rect 312170 10752 312176 10764
rect 312228 10752 312234 10804
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 29086 10724 29092 10736
rect 19392 10696 29092 10724
rect 19392 10684 19398 10696
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 33134 10684 33140 10736
rect 33192 10724 33198 10736
rect 42794 10724 42800 10736
rect 33192 10696 42800 10724
rect 33192 10684 33198 10696
rect 42794 10684 42800 10696
rect 42852 10684 42858 10736
rect 51718 10684 51724 10736
rect 51776 10724 51782 10736
rect 75914 10724 75920 10736
rect 51776 10696 75920 10724
rect 51776 10684 51782 10696
rect 75914 10684 75920 10696
rect 75972 10684 75978 10736
rect 82262 10684 82268 10736
rect 82320 10724 82326 10736
rect 249058 10724 249064 10736
rect 82320 10696 249064 10724
rect 82320 10684 82326 10696
rect 249058 10684 249064 10696
rect 249116 10684 249122 10736
rect 282914 10684 282920 10736
rect 282972 10724 282978 10736
rect 417418 10724 417424 10736
rect 282972 10696 417424 10724
rect 282972 10684 282978 10696
rect 417418 10684 417424 10696
rect 417476 10684 417482 10736
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 23474 10656 23480 10668
rect 14976 10628 23480 10656
rect 14976 10616 14982 10628
rect 23474 10616 23480 10628
rect 23532 10616 23538 10668
rect 30098 10616 30104 10668
rect 30156 10656 30162 10668
rect 44542 10656 44548 10668
rect 30156 10628 44548 10656
rect 30156 10616 30162 10628
rect 44542 10616 44548 10628
rect 44600 10616 44606 10668
rect 56134 10616 56140 10668
rect 56192 10656 56198 10668
rect 94498 10656 94504 10668
rect 56192 10628 94504 10656
rect 56192 10616 56198 10628
rect 94498 10616 94504 10628
rect 94556 10616 94562 10668
rect 95418 10616 95424 10668
rect 95476 10656 95482 10668
rect 96798 10656 96804 10668
rect 95476 10628 96804 10656
rect 95476 10616 95482 10628
rect 96798 10616 96804 10628
rect 96856 10616 96862 10668
rect 101674 10616 101680 10668
rect 101732 10656 101738 10668
rect 102318 10656 102324 10668
rect 101732 10628 102324 10656
rect 101732 10616 101738 10628
rect 102318 10616 102324 10628
rect 102376 10616 102382 10668
rect 104802 10616 104808 10668
rect 104860 10656 104866 10668
rect 109126 10656 109132 10668
rect 104860 10628 109132 10656
rect 104860 10616 104866 10628
rect 109126 10616 109132 10628
rect 109184 10616 109190 10668
rect 110414 10616 110420 10668
rect 110472 10656 110478 10668
rect 285674 10656 285680 10668
rect 110472 10628 285680 10656
rect 110472 10616 110478 10628
rect 285674 10616 285680 10628
rect 285732 10616 285738 10668
rect 299382 10616 299388 10668
rect 299440 10656 299446 10668
rect 309870 10656 309876 10668
rect 299440 10628 309876 10656
rect 299440 10616 299446 10628
rect 309870 10616 309876 10628
rect 309928 10616 309934 10668
rect 5442 10548 5448 10600
rect 5500 10588 5506 10600
rect 23566 10588 23572 10600
rect 5500 10560 23572 10588
rect 5500 10548 5506 10560
rect 23566 10548 23572 10560
rect 23624 10548 23630 10600
rect 40586 10548 40592 10600
rect 40644 10588 40650 10600
rect 65794 10588 65800 10600
rect 40644 10560 65800 10588
rect 40644 10548 40650 10560
rect 65794 10548 65800 10560
rect 65852 10548 65858 10600
rect 90082 10548 90088 10600
rect 90140 10588 90146 10600
rect 305546 10588 305552 10600
rect 90140 10560 305552 10588
rect 90140 10548 90146 10560
rect 305546 10548 305552 10560
rect 305604 10548 305610 10600
rect 14274 10480 14280 10532
rect 14332 10520 14338 10532
rect 41782 10520 41788 10532
rect 14332 10492 41788 10520
rect 14332 10480 14338 10492
rect 41782 10480 41788 10492
rect 41840 10480 41846 10532
rect 55766 10480 55772 10532
rect 55824 10520 55830 10532
rect 96614 10520 96620 10532
rect 55824 10492 96620 10520
rect 55824 10480 55830 10492
rect 96614 10480 96620 10492
rect 96672 10480 96678 10532
rect 96798 10480 96804 10532
rect 96856 10520 96862 10532
rect 103606 10520 103612 10532
rect 96856 10492 103612 10520
rect 96856 10480 96862 10492
rect 103606 10480 103612 10492
rect 103664 10480 103670 10532
rect 108298 10480 108304 10532
rect 108356 10520 108362 10532
rect 313274 10520 313280 10532
rect 108356 10492 313280 10520
rect 108356 10480 108362 10492
rect 313274 10480 313280 10492
rect 313332 10480 313338 10532
rect 335998 10480 336004 10532
rect 336056 10520 336062 10532
rect 362954 10520 362960 10532
rect 336056 10492 362960 10520
rect 336056 10480 336062 10492
rect 362954 10480 362960 10492
rect 363012 10480 363018 10532
rect 398926 10480 398932 10532
rect 398984 10520 398990 10532
rect 427170 10520 427176 10532
rect 398984 10492 427176 10520
rect 398984 10480 398990 10492
rect 427170 10480 427176 10492
rect 427228 10480 427234 10532
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 57882 10452 57888 10464
rect 11112 10424 57888 10452
rect 11112 10412 11118 10424
rect 57882 10412 57888 10424
rect 57940 10412 57946 10464
rect 61930 10412 61936 10464
rect 61988 10452 61994 10464
rect 68554 10452 68560 10464
rect 61988 10424 68560 10452
rect 61988 10412 61994 10424
rect 68554 10412 68560 10424
rect 68612 10412 68618 10464
rect 92290 10412 92296 10464
rect 92348 10452 92354 10464
rect 337010 10452 337016 10464
rect 92348 10424 337016 10452
rect 92348 10412 92354 10424
rect 337010 10412 337016 10424
rect 337068 10412 337074 10464
rect 354030 10412 354036 10464
rect 354088 10452 354094 10464
rect 367830 10452 367836 10464
rect 354088 10424 367836 10452
rect 354088 10412 354094 10424
rect 367830 10412 367836 10424
rect 367888 10412 367894 10464
rect 417234 10412 417240 10464
rect 417292 10452 417298 10464
rect 449158 10452 449164 10464
rect 417292 10424 449164 10452
rect 417292 10412 417298 10424
rect 449158 10412 449164 10424
rect 449216 10412 449222 10464
rect 13262 10344 13268 10396
rect 13320 10384 13326 10396
rect 59906 10384 59912 10396
rect 13320 10356 59912 10384
rect 13320 10344 13326 10356
rect 59906 10344 59912 10356
rect 59964 10344 59970 10396
rect 61470 10344 61476 10396
rect 61528 10384 61534 10396
rect 68646 10384 68652 10396
rect 61528 10356 68652 10384
rect 61528 10344 61534 10356
rect 68646 10344 68652 10356
rect 68704 10344 68710 10396
rect 68922 10344 68928 10396
rect 68980 10384 68986 10396
rect 82446 10384 82452 10396
rect 68980 10356 82452 10384
rect 68980 10344 68986 10356
rect 82446 10344 82452 10356
rect 82504 10344 82510 10396
rect 83550 10344 83556 10396
rect 83608 10384 83614 10396
rect 278038 10384 278044 10396
rect 83608 10356 278044 10384
rect 83608 10344 83614 10356
rect 278038 10344 278044 10356
rect 278096 10344 278102 10396
rect 285766 10344 285772 10396
rect 285824 10384 285830 10396
rect 548610 10384 548616 10396
rect 285824 10356 548616 10384
rect 285824 10344 285830 10356
rect 548610 10344 548616 10356
rect 548668 10344 548674 10396
rect 9582 10276 9588 10328
rect 9640 10316 9646 10328
rect 88334 10316 88340 10328
rect 9640 10288 88340 10316
rect 9640 10276 9646 10288
rect 88334 10276 88340 10288
rect 88392 10276 88398 10328
rect 94498 10276 94504 10328
rect 94556 10316 94562 10328
rect 96338 10316 96344 10328
rect 94556 10288 96344 10316
rect 94556 10276 94562 10288
rect 96338 10276 96344 10288
rect 96396 10276 96402 10328
rect 96614 10276 96620 10328
rect 96672 10316 96678 10328
rect 96890 10316 96896 10328
rect 96672 10288 96896 10316
rect 96672 10276 96678 10288
rect 96890 10276 96896 10288
rect 96948 10276 96954 10328
rect 98638 10276 98644 10328
rect 98696 10316 98702 10328
rect 108298 10316 108304 10328
rect 98696 10288 108304 10316
rect 98696 10276 98702 10288
rect 108298 10276 108304 10288
rect 108356 10276 108362 10328
rect 114554 10276 114560 10328
rect 114612 10316 114618 10328
rect 116118 10316 116124 10328
rect 114612 10288 116124 10316
rect 114612 10276 114618 10288
rect 116118 10276 116124 10288
rect 116176 10276 116182 10328
rect 132586 10276 132592 10328
rect 132644 10316 132650 10328
rect 534810 10316 534816 10328
rect 132644 10288 534816 10316
rect 132644 10276 132650 10288
rect 534810 10276 534816 10288
rect 534868 10276 534874 10328
rect 60918 10208 60924 10260
rect 60976 10248 60982 10260
rect 128446 10248 128452 10260
rect 60976 10220 128452 10248
rect 60976 10208 60982 10220
rect 128446 10208 128452 10220
rect 128504 10208 128510 10260
rect 147030 10208 147036 10260
rect 147088 10248 147094 10260
rect 154022 10248 154028 10260
rect 147088 10220 154028 10248
rect 147088 10208 147094 10220
rect 154022 10208 154028 10220
rect 154080 10208 154086 10260
rect 182266 10208 182272 10260
rect 182324 10248 182330 10260
rect 183738 10248 183744 10260
rect 182324 10220 183744 10248
rect 182324 10208 182330 10220
rect 183738 10208 183744 10220
rect 183796 10208 183802 10260
rect 52454 10140 52460 10192
rect 52512 10180 52518 10192
rect 78122 10180 78128 10192
rect 52512 10152 78128 10180
rect 52512 10140 52518 10152
rect 78122 10140 78128 10152
rect 78180 10140 78186 10192
rect 78582 10140 78588 10192
rect 78640 10180 78646 10192
rect 131114 10180 131120 10192
rect 78640 10152 131120 10180
rect 78640 10140 78646 10152
rect 131114 10140 131120 10152
rect 131172 10140 131178 10192
rect 92474 10112 92480 10124
rect 80026 10084 92480 10112
rect 54478 10004 54484 10056
rect 54536 10044 54542 10056
rect 80026 10044 80054 10084
rect 92474 10072 92480 10084
rect 92532 10072 92538 10124
rect 93762 10072 93768 10124
rect 93820 10112 93826 10124
rect 98086 10112 98092 10124
rect 93820 10084 98092 10112
rect 93820 10072 93826 10084
rect 98086 10072 98092 10084
rect 98144 10072 98150 10124
rect 135162 10112 135168 10124
rect 99346 10084 135168 10112
rect 99346 10044 99374 10084
rect 135162 10072 135168 10084
rect 135220 10072 135226 10124
rect 54536 10016 80054 10044
rect 89824 10016 99374 10044
rect 54536 10004 54542 10016
rect 64782 9936 64788 9988
rect 64840 9976 64846 9988
rect 68738 9976 68744 9988
rect 64840 9948 68744 9976
rect 64840 9936 64846 9948
rect 68738 9936 68744 9948
rect 68796 9936 68802 9988
rect 70394 9936 70400 9988
rect 70452 9976 70458 9988
rect 70452 9948 84884 9976
rect 70452 9936 70458 9948
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 81618 9908 81624 9920
rect 10836 9880 81624 9908
rect 10836 9868 10842 9880
rect 81618 9868 81624 9880
rect 81676 9868 81682 9920
rect 84856 9840 84884 9948
rect 88242 9868 88248 9920
rect 88300 9908 88306 9920
rect 89824 9908 89852 10016
rect 104802 10004 104808 10056
rect 104860 10044 104866 10056
rect 113082 10044 113088 10056
rect 104860 10016 113088 10044
rect 104860 10004 104866 10016
rect 113082 10004 113088 10016
rect 113140 10004 113146 10056
rect 128538 10004 128544 10056
rect 128596 10044 128602 10056
rect 140774 10044 140780 10056
rect 128596 10016 140780 10044
rect 128596 10004 128602 10016
rect 140774 10004 140780 10016
rect 140832 10004 140838 10056
rect 166074 9976 166080 9988
rect 88300 9880 89852 9908
rect 99346 9948 166080 9976
rect 88300 9868 88306 9880
rect 99346 9840 99374 9948
rect 166074 9936 166080 9948
rect 166132 9936 166138 9988
rect 84856 9812 99374 9840
rect 125134 9800 125140 9852
rect 125192 9840 125198 9852
rect 127526 9840 127532 9852
rect 125192 9812 127532 9840
rect 125192 9800 125198 9812
rect 127526 9800 127532 9812
rect 127584 9800 127590 9852
rect 156506 9732 156512 9784
rect 156564 9772 156570 9784
rect 180058 9772 180064 9784
rect 156564 9744 180064 9772
rect 156564 9732 156570 9744
rect 180058 9732 180064 9744
rect 180116 9732 180122 9784
rect 84562 9664 84568 9716
rect 84620 9704 84626 9716
rect 91002 9704 91008 9716
rect 84620 9676 91008 9704
rect 84620 9664 84626 9676
rect 91002 9664 91008 9676
rect 91060 9664 91066 9716
rect 123478 9704 123484 9716
rect 115952 9676 123484 9704
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 72418 9636 72424 9648
rect 12492 9608 72424 9636
rect 12492 9596 12498 9608
rect 72418 9596 72424 9608
rect 72476 9596 72482 9648
rect 86770 9596 86776 9648
rect 86828 9636 86834 9648
rect 91646 9636 91652 9648
rect 86828 9608 91652 9636
rect 86828 9596 86834 9608
rect 91646 9596 91652 9608
rect 91704 9596 91710 9648
rect 98270 9596 98276 9648
rect 98328 9636 98334 9648
rect 100386 9636 100392 9648
rect 98328 9608 100392 9636
rect 98328 9596 98334 9608
rect 100386 9596 100392 9608
rect 100444 9596 100450 9648
rect 101030 9596 101036 9648
rect 101088 9636 101094 9648
rect 111794 9636 111800 9648
rect 101088 9608 111800 9636
rect 101088 9596 101094 9608
rect 111794 9596 111800 9608
rect 111852 9596 111858 9648
rect 115842 9596 115848 9648
rect 115900 9636 115906 9648
rect 115952 9636 115980 9676
rect 123478 9664 123484 9676
rect 123536 9664 123542 9716
rect 131114 9664 131120 9716
rect 131172 9704 131178 9716
rect 240778 9704 240784 9716
rect 131172 9676 240784 9704
rect 131172 9664 131178 9676
rect 240778 9664 240784 9676
rect 240836 9664 240842 9716
rect 115900 9608 115980 9636
rect 115900 9596 115906 9608
rect 123754 9596 123760 9648
rect 123812 9636 123818 9648
rect 124582 9636 124588 9648
rect 123812 9608 124588 9636
rect 123812 9596 123818 9608
rect 124582 9596 124588 9608
rect 124640 9596 124646 9648
rect 143074 9596 143080 9648
rect 143132 9636 143138 9648
rect 143902 9636 143908 9648
rect 143132 9608 143908 9636
rect 143132 9596 143138 9608
rect 143902 9596 143908 9608
rect 143960 9596 143966 9648
rect 156966 9596 156972 9648
rect 157024 9636 157030 9648
rect 159358 9636 159364 9648
rect 157024 9608 159364 9636
rect 157024 9596 157030 9608
rect 159358 9596 159364 9608
rect 159416 9596 159422 9648
rect 183462 9596 183468 9648
rect 183520 9636 183526 9648
rect 232038 9636 232044 9648
rect 183520 9608 232044 9636
rect 183520 9596 183526 9608
rect 232038 9596 232044 9608
rect 232096 9596 232102 9648
rect 356790 9596 356796 9648
rect 356848 9636 356854 9648
rect 360102 9636 360108 9648
rect 356848 9608 360108 9636
rect 356848 9596 356854 9608
rect 360102 9596 360108 9608
rect 360160 9596 360166 9648
rect 367738 9596 367744 9648
rect 367796 9636 367802 9648
rect 372890 9636 372896 9648
rect 367796 9608 372896 9636
rect 367796 9596 367802 9608
rect 372890 9596 372896 9608
rect 372948 9596 372954 9648
rect 387794 9596 387800 9648
rect 387852 9636 387858 9648
rect 391842 9636 391848 9648
rect 387852 9608 391848 9636
rect 387852 9596 387858 9608
rect 391842 9596 391848 9608
rect 391900 9596 391906 9648
rect 403618 9596 403624 9648
rect 403676 9636 403682 9648
rect 406010 9636 406016 9648
rect 403676 9608 406016 9636
rect 403676 9596 403682 9608
rect 406010 9596 406016 9608
rect 406068 9596 406074 9648
rect 434898 9596 434904 9648
rect 434956 9636 434962 9648
rect 438762 9636 438768 9648
rect 434956 9608 438768 9636
rect 434956 9596 434962 9608
rect 438762 9596 438768 9608
rect 438820 9596 438826 9648
rect 502978 9596 502984 9648
rect 503036 9636 503042 9648
rect 506474 9636 506480 9648
rect 503036 9608 506480 9636
rect 503036 9596 503042 9608
rect 506474 9596 506480 9608
rect 506532 9596 506538 9648
rect 23658 9528 23664 9580
rect 23716 9568 23722 9580
rect 68922 9568 68928 9580
rect 23716 9540 68928 9568
rect 23716 9528 23722 9540
rect 68922 9528 68928 9540
rect 68980 9528 68986 9580
rect 90192 9540 90404 9568
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 70670 9500 70676 9512
rect 18840 9472 70676 9500
rect 18840 9460 18846 9472
rect 70670 9460 70676 9472
rect 70728 9460 70734 9512
rect 80882 9460 80888 9512
rect 80940 9500 80946 9512
rect 90192 9500 90220 9540
rect 80940 9472 90220 9500
rect 90376 9500 90404 9540
rect 91002 9528 91008 9580
rect 91060 9568 91066 9580
rect 102134 9568 102140 9580
rect 91060 9540 102140 9568
rect 91060 9528 91066 9540
rect 102134 9528 102140 9540
rect 102192 9528 102198 9580
rect 107746 9528 107752 9580
rect 107804 9568 107810 9580
rect 111518 9568 111524 9580
rect 107804 9540 111524 9568
rect 107804 9528 107810 9540
rect 111518 9528 111524 9540
rect 111576 9528 111582 9580
rect 112162 9528 112168 9580
rect 112220 9568 112226 9580
rect 114646 9568 114652 9580
rect 112220 9540 114652 9568
rect 112220 9528 112226 9540
rect 114646 9528 114652 9540
rect 114704 9528 114710 9580
rect 154298 9528 154304 9580
rect 154356 9568 154362 9580
rect 158070 9568 158076 9580
rect 154356 9540 158076 9568
rect 154356 9528 154362 9540
rect 158070 9528 158076 9540
rect 158128 9528 158134 9580
rect 209682 9528 209688 9580
rect 209740 9568 209746 9580
rect 210970 9568 210976 9580
rect 209740 9540 210976 9568
rect 209740 9528 209746 9540
rect 210970 9528 210976 9540
rect 211028 9528 211034 9580
rect 223390 9528 223396 9580
rect 223448 9568 223454 9580
rect 292206 9568 292212 9580
rect 223448 9540 292212 9568
rect 223448 9528 223454 9540
rect 292206 9528 292212 9540
rect 292264 9528 292270 9580
rect 356698 9528 356704 9580
rect 356756 9568 356762 9580
rect 360010 9568 360016 9580
rect 356756 9540 360016 9568
rect 356756 9528 356762 9540
rect 360010 9528 360016 9540
rect 360068 9528 360074 9580
rect 405826 9528 405832 9580
rect 405884 9568 405890 9580
rect 408678 9568 408684 9580
rect 405884 9540 408684 9568
rect 405884 9528 405890 9540
rect 408678 9528 408684 9540
rect 408736 9528 408742 9580
rect 234522 9500 234528 9512
rect 90376 9472 234528 9500
rect 80940 9460 80946 9472
rect 234522 9460 234528 9472
rect 234580 9460 234586 9512
rect 235994 9460 236000 9512
rect 236052 9500 236058 9512
rect 242986 9500 242992 9512
rect 236052 9472 242992 9500
rect 236052 9460 236058 9472
rect 242986 9460 242992 9472
rect 243044 9460 243050 9512
rect 463142 9460 463148 9512
rect 463200 9500 463206 9512
rect 467650 9500 467656 9512
rect 463200 9472 467656 9500
rect 463200 9460 463206 9472
rect 467650 9460 467656 9472
rect 467708 9460 467714 9512
rect 18598 9392 18604 9444
rect 18656 9432 18662 9444
rect 90174 9432 90180 9444
rect 18656 9404 90180 9432
rect 18656 9392 18662 9404
rect 90174 9392 90180 9404
rect 90232 9392 90238 9444
rect 91830 9392 91836 9444
rect 91888 9432 91894 9444
rect 282822 9432 282828 9444
rect 91888 9404 282828 9432
rect 91888 9392 91894 9404
rect 282822 9392 282828 9404
rect 282880 9392 282886 9444
rect 284294 9392 284300 9444
rect 284352 9432 284358 9444
rect 343358 9432 343364 9444
rect 284352 9404 343364 9432
rect 284352 9392 284358 9404
rect 343358 9392 343364 9404
rect 343416 9392 343422 9444
rect 510246 9392 510252 9444
rect 510304 9432 510310 9444
rect 517146 9432 517152 9444
rect 510304 9404 517152 9432
rect 510304 9392 510310 9404
rect 517146 9392 517152 9404
rect 517204 9392 517210 9444
rect 52822 9324 52828 9376
rect 52880 9364 52886 9376
rect 83274 9364 83280 9376
rect 52880 9336 83280 9364
rect 52880 9324 52886 9336
rect 83274 9324 83280 9336
rect 83332 9324 83338 9376
rect 86494 9324 86500 9376
rect 86552 9364 86558 9376
rect 277394 9364 277400 9376
rect 86552 9336 277400 9364
rect 86552 9324 86558 9336
rect 277394 9324 277400 9336
rect 277452 9324 277458 9376
rect 285674 9324 285680 9376
rect 285732 9364 285738 9376
rect 354030 9364 354036 9376
rect 285732 9336 354036 9364
rect 285732 9324 285738 9336
rect 354030 9324 354036 9336
rect 354088 9324 354094 9376
rect 438118 9324 438124 9376
rect 438176 9364 438182 9376
rect 449434 9364 449440 9376
rect 438176 9336 449440 9364
rect 438176 9324 438182 9336
rect 449434 9324 449440 9336
rect 449492 9324 449498 9376
rect 491202 9324 491208 9376
rect 491260 9364 491266 9376
rect 510062 9364 510068 9376
rect 491260 9336 510068 9364
rect 491260 9324 491266 9336
rect 510062 9324 510068 9336
rect 510120 9324 510126 9376
rect 17126 9256 17132 9308
rect 17184 9296 17190 9308
rect 26326 9296 26332 9308
rect 17184 9268 26332 9296
rect 17184 9256 17190 9268
rect 26326 9256 26332 9268
rect 26384 9256 26390 9308
rect 94774 9256 94780 9308
rect 94832 9296 94838 9308
rect 291746 9296 291752 9308
rect 94832 9268 291752 9296
rect 94832 9256 94838 9268
rect 291746 9256 291752 9268
rect 291804 9256 291810 9308
rect 404262 9256 404268 9308
rect 404320 9296 404326 9308
rect 427722 9296 427728 9308
rect 404320 9268 427728 9296
rect 404320 9256 404326 9268
rect 427722 9256 427728 9268
rect 427780 9256 427786 9308
rect 440234 9256 440240 9308
rect 440292 9296 440298 9308
rect 452746 9296 452752 9308
rect 440292 9268 452752 9296
rect 440292 9256 440298 9268
rect 452746 9256 452752 9268
rect 452804 9256 452810 9308
rect 456058 9256 456064 9308
rect 456116 9296 456122 9308
rect 471974 9296 471980 9308
rect 456116 9268 471980 9296
rect 456116 9256 456122 9268
rect 471974 9256 471980 9268
rect 472032 9256 472038 9308
rect 473998 9256 474004 9308
rect 474056 9296 474062 9308
rect 491294 9296 491300 9308
rect 474056 9268 491300 9296
rect 474056 9256 474062 9268
rect 491294 9256 491300 9268
rect 491352 9256 491358 9308
rect 507118 9256 507124 9308
rect 507176 9296 507182 9308
rect 534902 9296 534908 9308
rect 507176 9268 534908 9296
rect 507176 9256 507182 9268
rect 534902 9256 534908 9268
rect 534960 9256 534966 9308
rect 20254 9188 20260 9240
rect 20312 9228 20318 9240
rect 56594 9228 56600 9240
rect 20312 9200 56600 9228
rect 20312 9188 20318 9200
rect 56594 9188 56600 9200
rect 56652 9188 56658 9240
rect 65610 9188 65616 9240
rect 65668 9228 65674 9240
rect 84746 9228 84752 9240
rect 65668 9200 84752 9228
rect 65668 9188 65674 9200
rect 84746 9188 84752 9200
rect 84804 9188 84810 9240
rect 87966 9188 87972 9240
rect 88024 9228 88030 9240
rect 287790 9228 287796 9240
rect 88024 9200 287796 9228
rect 88024 9188 88030 9200
rect 287790 9188 287796 9200
rect 287848 9188 287854 9240
rect 313274 9188 313280 9240
rect 313332 9228 313338 9240
rect 377674 9228 377680 9240
rect 313332 9200 377680 9228
rect 313332 9188 313338 9200
rect 377674 9188 377680 9200
rect 377732 9188 377738 9240
rect 390922 9188 390928 9240
rect 390980 9228 390986 9240
rect 400122 9228 400128 9240
rect 390980 9200 400128 9228
rect 390980 9188 390986 9200
rect 400122 9188 400128 9200
rect 400180 9188 400186 9240
rect 408494 9188 408500 9240
rect 408552 9228 408558 9240
rect 435450 9228 435456 9240
rect 408552 9200 435456 9228
rect 408552 9188 408558 9200
rect 435450 9188 435456 9200
rect 435508 9188 435514 9240
rect 435910 9188 435916 9240
rect 435968 9228 435974 9240
rect 458082 9228 458088 9240
rect 435968 9200 458088 9228
rect 435968 9188 435974 9200
rect 458082 9188 458088 9200
rect 458140 9188 458146 9240
rect 458818 9188 458824 9240
rect 458876 9228 458882 9240
rect 470686 9228 470692 9240
rect 458876 9200 470692 9228
rect 458876 9188 458882 9200
rect 470686 9188 470692 9200
rect 470744 9188 470750 9240
rect 491938 9188 491944 9240
rect 491996 9228 492002 9240
rect 528554 9228 528560 9240
rect 491996 9200 528560 9228
rect 491996 9188 492002 9200
rect 528554 9188 528560 9200
rect 528612 9188 528618 9240
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 40770 9160 40776 9172
rect 13596 9132 40776 9160
rect 13596 9120 13602 9132
rect 40770 9120 40776 9132
rect 40828 9120 40834 9172
rect 55030 9120 55036 9172
rect 55088 9160 55094 9172
rect 93854 9160 93860 9172
rect 55088 9132 93860 9160
rect 55088 9120 55094 9132
rect 93854 9120 93860 9132
rect 93912 9120 93918 9172
rect 97994 9120 98000 9172
rect 98052 9160 98058 9172
rect 106274 9160 106280 9172
rect 98052 9132 106280 9160
rect 98052 9120 98058 9132
rect 106274 9120 106280 9132
rect 106332 9120 106338 9172
rect 109126 9120 109132 9172
rect 109184 9160 109190 9172
rect 318702 9160 318708 9172
rect 109184 9132 318708 9160
rect 109184 9120 109190 9132
rect 318702 9120 318708 9132
rect 318760 9120 318766 9172
rect 348510 9120 348516 9172
rect 348568 9160 348574 9172
rect 357526 9160 357532 9172
rect 348568 9132 357532 9160
rect 348568 9120 348574 9132
rect 357526 9120 357532 9132
rect 357584 9120 357590 9172
rect 380986 9120 380992 9172
rect 381044 9160 381050 9172
rect 412634 9160 412640 9172
rect 381044 9132 412640 9160
rect 381044 9120 381050 9132
rect 412634 9120 412640 9132
rect 412692 9120 412698 9172
rect 424962 9120 424968 9172
rect 425020 9160 425026 9172
rect 436002 9160 436008 9172
rect 425020 9132 436008 9160
rect 425020 9120 425026 9132
rect 436002 9120 436008 9132
rect 436060 9120 436066 9172
rect 448698 9120 448704 9172
rect 448756 9160 448762 9172
rect 476022 9160 476028 9172
rect 448756 9132 476028 9160
rect 448756 9120 448762 9132
rect 476022 9120 476028 9132
rect 476080 9120 476086 9172
rect 488534 9120 488540 9172
rect 488592 9160 488598 9172
rect 526254 9160 526260 9172
rect 488592 9132 526260 9160
rect 488592 9120 488598 9132
rect 526254 9120 526260 9132
rect 526312 9120 526318 9172
rect 531222 9120 531228 9172
rect 531280 9160 531286 9172
rect 541986 9160 541992 9172
rect 531280 9132 541992 9160
rect 531280 9120 531286 9132
rect 541986 9120 541992 9132
rect 542044 9120 542050 9172
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 67910 9092 67916 9104
rect 19668 9064 67916 9092
rect 19668 9052 19674 9064
rect 67910 9052 67916 9064
rect 67968 9052 67974 9104
rect 68830 9052 68836 9104
rect 68888 9092 68894 9104
rect 86954 9092 86960 9104
rect 68888 9064 86960 9092
rect 68888 9052 68894 9064
rect 86954 9052 86960 9064
rect 87012 9052 87018 9104
rect 88334 9052 88340 9104
rect 88392 9092 88398 9104
rect 88392 9064 99374 9092
rect 88392 9052 88398 9064
rect 20530 8984 20536 9036
rect 20588 9024 20594 9036
rect 71774 9024 71780 9036
rect 20588 8996 71780 9024
rect 20588 8984 20594 8996
rect 71774 8984 71780 8996
rect 71832 8984 71838 9036
rect 81526 8984 81532 9036
rect 81584 9024 81590 9036
rect 81584 8996 91140 9024
rect 81584 8984 81590 8996
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 20622 8956 20628 8968
rect 15252 8928 20628 8956
rect 15252 8916 15258 8928
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 21082 8916 21088 8968
rect 21140 8956 21146 8968
rect 82078 8956 82084 8968
rect 21140 8928 82084 8956
rect 21140 8916 21146 8928
rect 82078 8916 82084 8928
rect 82136 8916 82142 8968
rect 85206 8916 85212 8968
rect 85264 8956 85270 8968
rect 91002 8956 91008 8968
rect 85264 8928 91008 8956
rect 85264 8916 85270 8928
rect 91002 8916 91008 8928
rect 91060 8916 91066 8968
rect 91112 8956 91140 8996
rect 95234 8984 95240 9036
rect 95292 9024 95298 9036
rect 97718 9024 97724 9036
rect 95292 8996 97724 9024
rect 95292 8984 95298 8996
rect 97718 8984 97724 8996
rect 97776 8984 97782 9036
rect 99346 9024 99374 9064
rect 100754 9052 100760 9104
rect 100812 9092 100818 9104
rect 350442 9092 350448 9104
rect 100812 9064 350448 9092
rect 100812 9052 100818 9064
rect 350442 9052 350448 9064
rect 350500 9052 350506 9104
rect 378042 9052 378048 9104
rect 378100 9092 378106 9104
rect 393038 9092 393044 9104
rect 378100 9064 393044 9092
rect 378100 9052 378106 9064
rect 393038 9052 393044 9064
rect 393096 9052 393102 9104
rect 394970 9052 394976 9104
rect 395028 9092 395034 9104
rect 403158 9092 403164 9104
rect 395028 9064 403164 9092
rect 395028 9052 395034 9064
rect 403158 9052 403164 9064
rect 403216 9052 403222 9104
rect 413554 9052 413560 9104
rect 413612 9092 413618 9104
rect 449802 9092 449808 9104
rect 413612 9064 449808 9092
rect 413612 9052 413618 9064
rect 449802 9052 449808 9064
rect 449860 9052 449866 9104
rect 449894 9052 449900 9104
rect 449952 9092 449958 9104
rect 498194 9092 498200 9104
rect 449952 9064 498200 9092
rect 449952 9052 449958 9064
rect 498194 9052 498200 9064
rect 498252 9052 498258 9104
rect 498286 9052 498292 9104
rect 498344 9092 498350 9104
rect 531314 9092 531320 9104
rect 498344 9064 531320 9092
rect 498344 9052 498350 9064
rect 531314 9052 531320 9064
rect 531372 9052 531378 9104
rect 534718 9052 534724 9104
rect 534776 9092 534782 9104
rect 571242 9092 571248 9104
rect 534776 9064 571248 9092
rect 534776 9052 534782 9064
rect 571242 9052 571248 9064
rect 571300 9052 571306 9104
rect 103514 9024 103520 9036
rect 99346 8996 103520 9024
rect 103514 8984 103520 8996
rect 103572 8984 103578 9036
rect 107562 8984 107568 9036
rect 107620 9024 107626 9036
rect 355226 9024 355232 9036
rect 107620 8996 355232 9024
rect 107620 8984 107626 8996
rect 355226 8984 355232 8996
rect 355284 8984 355290 9036
rect 377950 8984 377956 9036
rect 378008 9024 378014 9036
rect 430574 9024 430580 9036
rect 378008 8996 430580 9024
rect 378008 8984 378014 8996
rect 430574 8984 430580 8996
rect 430632 8984 430638 9036
rect 431310 8984 431316 9036
rect 431368 9024 431374 9036
rect 445018 9024 445024 9036
rect 431368 8996 445024 9024
rect 431368 8984 431374 8996
rect 445018 8984 445024 8996
rect 445076 8984 445082 9036
rect 445662 8984 445668 9036
rect 445720 9024 445726 9036
rect 478874 9024 478880 9036
rect 445720 8996 478880 9024
rect 445720 8984 445726 8996
rect 478874 8984 478880 8996
rect 478932 8984 478938 9036
rect 493962 8984 493968 9036
rect 494020 9024 494026 9036
rect 565814 9024 565820 9036
rect 494020 8996 565820 9024
rect 494020 8984 494026 8996
rect 565814 8984 565820 8996
rect 565872 8984 565878 9036
rect 101214 8956 101220 8968
rect 91112 8928 101220 8956
rect 101214 8916 101220 8928
rect 101272 8916 101278 8968
rect 101582 8916 101588 8968
rect 101640 8956 101646 8968
rect 382366 8956 382372 8968
rect 101640 8928 382372 8956
rect 101640 8916 101646 8928
rect 382366 8916 382372 8928
rect 382424 8916 382430 8968
rect 385310 8916 385316 8968
rect 385368 8956 385374 8968
rect 394694 8956 394700 8968
rect 385368 8928 394700 8956
rect 385368 8916 385374 8928
rect 394694 8916 394700 8928
rect 394752 8916 394758 8968
rect 398834 8916 398840 8968
rect 398892 8956 398898 8968
rect 416866 8956 416872 8968
rect 398892 8928 416872 8956
rect 398892 8916 398898 8928
rect 416866 8916 416872 8928
rect 416924 8916 416930 8968
rect 426986 8916 426992 8968
rect 427044 8956 427050 8968
rect 503622 8956 503628 8968
rect 427044 8928 503628 8956
rect 427044 8916 427050 8928
rect 503622 8916 503628 8928
rect 503680 8916 503686 8968
rect 516134 8916 516140 8968
rect 516192 8956 516198 8968
rect 577406 8956 577412 8968
rect 516192 8928 577412 8956
rect 516192 8916 516198 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 49878 8848 49884 8900
rect 49936 8888 49942 8900
rect 64322 8888 64328 8900
rect 49936 8860 64328 8888
rect 49936 8848 49942 8860
rect 64322 8848 64328 8860
rect 64380 8848 64386 8900
rect 70486 8848 70492 8900
rect 70544 8888 70550 8900
rect 154206 8888 154212 8900
rect 70544 8860 89714 8888
rect 70544 8848 70550 8860
rect 56686 8780 56692 8832
rect 56744 8820 56750 8832
rect 56744 8792 80054 8820
rect 56744 8780 56750 8792
rect 80026 8684 80054 8792
rect 83366 8780 83372 8832
rect 83424 8820 83430 8832
rect 84654 8820 84660 8832
rect 83424 8792 84660 8820
rect 83424 8780 83430 8792
rect 84654 8780 84660 8792
rect 84712 8780 84718 8832
rect 89686 8820 89714 8860
rect 91112 8860 154212 8888
rect 91112 8820 91140 8860
rect 154206 8848 154212 8860
rect 154264 8848 154270 8900
rect 160186 8848 160192 8900
rect 160244 8888 160250 8900
rect 186866 8888 186872 8900
rect 160244 8860 186872 8888
rect 160244 8848 160250 8860
rect 186866 8848 186872 8860
rect 186924 8848 186930 8900
rect 89686 8792 91140 8820
rect 135162 8780 135168 8832
rect 135220 8820 135226 8832
rect 139302 8820 139308 8832
rect 135220 8792 139308 8820
rect 135220 8780 135226 8792
rect 139302 8780 139308 8792
rect 139360 8780 139366 8832
rect 82722 8712 82728 8764
rect 82780 8752 82786 8764
rect 101306 8752 101312 8764
rect 82780 8724 101312 8752
rect 82780 8712 82786 8724
rect 101306 8712 101312 8724
rect 101364 8712 101370 8764
rect 88426 8684 88432 8696
rect 80026 8656 88432 8684
rect 88426 8644 88432 8656
rect 88484 8644 88490 8696
rect 91002 8644 91008 8696
rect 91060 8684 91066 8696
rect 94498 8684 94504 8696
rect 91060 8656 94504 8684
rect 91060 8644 91066 8656
rect 94498 8644 94504 8656
rect 94556 8644 94562 8696
rect 96614 8644 96620 8696
rect 96672 8684 96678 8696
rect 100938 8684 100944 8696
rect 96672 8656 100944 8684
rect 96672 8644 96678 8656
rect 100938 8644 100944 8656
rect 100996 8644 101002 8696
rect 128446 8644 128452 8696
rect 128504 8684 128510 8696
rect 131206 8684 131212 8696
rect 128504 8656 131212 8684
rect 128504 8644 128510 8656
rect 131206 8644 131212 8656
rect 131264 8644 131270 8696
rect 351914 8644 351920 8696
rect 351972 8684 351978 8696
rect 354674 8684 354680 8696
rect 351972 8656 354680 8684
rect 351972 8644 351978 8656
rect 354674 8644 354680 8656
rect 354732 8644 354738 8696
rect 68278 8576 68284 8628
rect 68336 8616 68342 8628
rect 162854 8616 162860 8628
rect 68336 8588 162860 8616
rect 68336 8576 68342 8588
rect 162854 8576 162860 8588
rect 162912 8576 162918 8628
rect 68094 8508 68100 8560
rect 68152 8548 68158 8560
rect 172514 8548 172520 8560
rect 68152 8520 172520 8548
rect 68152 8508 68158 8520
rect 172514 8508 172520 8520
rect 172572 8508 172578 8560
rect 59906 8440 59912 8492
rect 59964 8480 59970 8492
rect 95326 8480 95332 8492
rect 59964 8452 95332 8480
rect 59964 8440 59970 8452
rect 95326 8440 95332 8452
rect 95384 8440 95390 8492
rect 444650 8372 444656 8424
rect 444708 8412 444714 8424
rect 452654 8412 452660 8424
rect 444708 8384 452660 8412
rect 444708 8372 444714 8384
rect 452654 8372 452660 8384
rect 452712 8372 452718 8424
rect 78306 8304 78312 8356
rect 78364 8344 78370 8356
rect 84378 8344 84384 8356
rect 78364 8316 84384 8344
rect 78364 8304 78370 8316
rect 84378 8304 84384 8316
rect 84436 8304 84442 8356
rect 102134 8304 102140 8356
rect 102192 8344 102198 8356
rect 107470 8344 107476 8356
rect 102192 8316 107476 8344
rect 102192 8304 102198 8316
rect 107470 8304 107476 8316
rect 107528 8304 107534 8356
rect 114646 8344 114652 8356
rect 110432 8316 114652 8344
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 94590 8276 94596 8288
rect 8996 8248 94596 8276
rect 8996 8236 9002 8248
rect 94590 8236 94596 8248
rect 94648 8236 94654 8288
rect 96062 8236 96068 8288
rect 96120 8276 96126 8288
rect 97442 8276 97448 8288
rect 96120 8248 97448 8276
rect 96120 8236 96126 8248
rect 97442 8236 97448 8248
rect 97500 8236 97506 8288
rect 98086 8236 98092 8288
rect 98144 8276 98150 8288
rect 102594 8276 102600 8288
rect 98144 8248 102600 8276
rect 98144 8236 98150 8248
rect 102594 8236 102600 8248
rect 102652 8236 102658 8288
rect 102686 8236 102692 8288
rect 102744 8276 102750 8288
rect 110432 8276 110460 8316
rect 114646 8304 114652 8316
rect 114704 8304 114710 8356
rect 125042 8344 125048 8356
rect 117240 8316 125048 8344
rect 102744 8248 110460 8276
rect 102744 8236 102750 8248
rect 115750 8236 115756 8288
rect 115808 8276 115814 8288
rect 117240 8276 117268 8316
rect 125042 8304 125048 8316
rect 125100 8304 125106 8356
rect 184750 8344 184756 8356
rect 126532 8316 128400 8344
rect 115808 8248 117268 8276
rect 115808 8236 115814 8248
rect 119338 8236 119344 8288
rect 119396 8276 119402 8288
rect 123018 8276 123024 8288
rect 119396 8248 123024 8276
rect 119396 8236 119402 8248
rect 123018 8236 123024 8248
rect 123076 8236 123082 8288
rect 65794 8168 65800 8220
rect 65852 8208 65858 8220
rect 71038 8208 71044 8220
rect 65852 8180 71044 8208
rect 65852 8168 65858 8180
rect 71038 8168 71044 8180
rect 71096 8168 71102 8220
rect 81342 8168 81348 8220
rect 81400 8208 81406 8220
rect 85022 8208 85028 8220
rect 81400 8180 85028 8208
rect 81400 8168 81406 8180
rect 85022 8168 85028 8180
rect 85080 8168 85086 8220
rect 116026 8168 116032 8220
rect 116084 8208 116090 8220
rect 119890 8208 119896 8220
rect 116084 8180 119896 8208
rect 116084 8168 116090 8180
rect 119890 8168 119896 8180
rect 119948 8168 119954 8220
rect 122466 8168 122472 8220
rect 122524 8208 122530 8220
rect 126532 8208 126560 8316
rect 128372 8276 128400 8316
rect 142126 8316 184756 8344
rect 130286 8276 130292 8288
rect 128372 8248 130292 8276
rect 130286 8236 130292 8248
rect 130344 8236 130350 8288
rect 137922 8236 137928 8288
rect 137980 8276 137986 8288
rect 142126 8276 142154 8316
rect 184750 8304 184756 8316
rect 184808 8304 184814 8356
rect 191742 8304 191748 8356
rect 191800 8344 191806 8356
rect 213822 8344 213828 8356
rect 191800 8316 213828 8344
rect 191800 8304 191806 8316
rect 213822 8304 213828 8316
rect 213880 8304 213886 8356
rect 137980 8248 142154 8276
rect 137980 8236 137986 8248
rect 146938 8236 146944 8288
rect 146996 8276 147002 8288
rect 149606 8276 149612 8288
rect 146996 8248 149612 8276
rect 146996 8236 147002 8248
rect 149606 8236 149612 8248
rect 149664 8236 149670 8288
rect 327534 8236 327540 8288
rect 327592 8276 327598 8288
rect 330846 8276 330852 8288
rect 327592 8248 330852 8276
rect 327592 8236 327598 8248
rect 330846 8236 330852 8248
rect 330904 8236 330910 8288
rect 122524 8180 126560 8208
rect 122524 8168 122530 8180
rect 149238 8168 149244 8220
rect 149296 8208 149302 8220
rect 151262 8208 151268 8220
rect 149296 8180 151268 8208
rect 149296 8168 149302 8180
rect 151262 8168 151268 8180
rect 151320 8168 151326 8220
rect 80606 8100 80612 8152
rect 80664 8140 80670 8152
rect 155310 8140 155316 8152
rect 80664 8112 155316 8140
rect 80664 8100 80670 8112
rect 155310 8100 155316 8112
rect 155368 8100 155374 8152
rect 202230 8100 202236 8152
rect 202288 8140 202294 8152
rect 223482 8140 223488 8152
rect 202288 8112 223488 8140
rect 202288 8100 202294 8112
rect 223482 8100 223488 8112
rect 223540 8100 223546 8152
rect 94038 8032 94044 8084
rect 94096 8072 94102 8084
rect 207658 8072 207664 8084
rect 94096 8044 207664 8072
rect 94096 8032 94102 8044
rect 207658 8032 207664 8044
rect 207716 8032 207722 8084
rect 22186 7964 22192 8016
rect 22244 8004 22250 8016
rect 90358 8004 90364 8016
rect 22244 7976 90364 8004
rect 22244 7964 22250 7976
rect 90358 7964 90364 7976
rect 90416 7964 90422 8016
rect 94498 7964 94504 8016
rect 94556 8004 94562 8016
rect 213730 8004 213736 8016
rect 94556 7976 213736 8004
rect 94556 7964 94562 7976
rect 213730 7964 213736 7976
rect 213788 7964 213794 8016
rect 37182 7896 37188 7948
rect 37240 7936 37246 7948
rect 70670 7936 70676 7948
rect 37240 7908 70676 7936
rect 37240 7896 37246 7908
rect 70670 7896 70676 7908
rect 70728 7896 70734 7948
rect 74718 7896 74724 7948
rect 74776 7936 74782 7948
rect 204162 7936 204168 7948
rect 74776 7908 204168 7936
rect 74776 7896 74782 7908
rect 204162 7896 204168 7908
rect 204220 7896 204226 7948
rect 213822 7896 213828 7948
rect 213880 7936 213886 7948
rect 236362 7936 236368 7948
rect 213880 7908 236368 7936
rect 213880 7896 213886 7908
rect 236362 7896 236368 7908
rect 236420 7896 236426 7948
rect 318610 7896 318616 7948
rect 318668 7936 318674 7948
rect 332686 7936 332692 7948
rect 318668 7908 332692 7936
rect 318668 7896 318674 7908
rect 332686 7896 332692 7908
rect 332744 7896 332750 7948
rect 29086 7828 29092 7880
rect 29144 7868 29150 7880
rect 92750 7868 92756 7880
rect 29144 7840 92756 7868
rect 29144 7828 29150 7840
rect 92750 7828 92756 7840
rect 92808 7828 92814 7880
rect 125594 7828 125600 7880
rect 125652 7868 125658 7880
rect 127802 7868 127808 7880
rect 125652 7840 127808 7868
rect 125652 7828 125658 7840
rect 127802 7828 127808 7840
rect 127860 7828 127866 7880
rect 129734 7828 129740 7880
rect 129792 7868 129798 7880
rect 265618 7868 265624 7880
rect 129792 7840 265624 7868
rect 129792 7828 129798 7840
rect 265618 7828 265624 7840
rect 265676 7828 265682 7880
rect 318702 7828 318708 7880
rect 318760 7868 318766 7880
rect 342070 7868 342076 7880
rect 318760 7840 342076 7868
rect 318760 7828 318766 7840
rect 342070 7828 342076 7840
rect 342128 7828 342134 7880
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 43162 7800 43168 7812
rect 24268 7772 43168 7800
rect 24268 7760 24274 7772
rect 43162 7760 43168 7772
rect 43220 7760 43226 7812
rect 54294 7760 54300 7812
rect 54352 7800 54358 7812
rect 90174 7800 90180 7812
rect 54352 7772 90180 7800
rect 54352 7760 54358 7772
rect 90174 7760 90180 7772
rect 90232 7760 90238 7812
rect 90634 7760 90640 7812
rect 90692 7800 90698 7812
rect 319714 7800 319720 7812
rect 90692 7772 319720 7800
rect 90692 7760 90698 7772
rect 319714 7760 319720 7772
rect 319772 7760 319778 7812
rect 362954 7760 362960 7812
rect 363012 7800 363018 7812
rect 389082 7800 389088 7812
rect 363012 7772 389088 7800
rect 363012 7760 363018 7772
rect 389082 7760 389088 7772
rect 389140 7760 389146 7812
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 40494 7732 40500 7744
rect 4212 7704 40500 7732
rect 4212 7692 4218 7704
rect 40494 7692 40500 7704
rect 40552 7692 40558 7744
rect 42794 7692 42800 7744
rect 42852 7732 42858 7744
rect 64874 7732 64880 7744
rect 42852 7704 64880 7732
rect 42852 7692 42858 7704
rect 64874 7692 64880 7704
rect 64932 7692 64938 7744
rect 90266 7692 90272 7744
rect 90324 7732 90330 7744
rect 321462 7732 321468 7744
rect 90324 7704 321468 7732
rect 90324 7692 90330 7704
rect 321462 7692 321468 7704
rect 321520 7692 321526 7744
rect 345842 7692 345848 7744
rect 345900 7732 345906 7744
rect 383562 7732 383568 7744
rect 345900 7704 383568 7732
rect 345900 7692 345906 7704
rect 383562 7692 383568 7704
rect 383620 7692 383626 7744
rect 15102 7624 15108 7676
rect 15160 7664 15166 7676
rect 35894 7664 35900 7676
rect 15160 7636 35900 7664
rect 15160 7624 15166 7636
rect 35894 7624 35900 7636
rect 35952 7624 35958 7676
rect 36814 7624 36820 7676
rect 36872 7664 36878 7676
rect 81342 7664 81348 7676
rect 36872 7636 81348 7664
rect 36872 7624 36878 7636
rect 81342 7624 81348 7636
rect 81400 7624 81406 7676
rect 88702 7624 88708 7676
rect 88760 7664 88766 7676
rect 94498 7664 94504 7676
rect 88760 7636 94504 7664
rect 88760 7624 88766 7636
rect 94498 7624 94504 7636
rect 94556 7624 94562 7676
rect 96706 7624 96712 7676
rect 96764 7664 96770 7676
rect 364610 7664 364616 7676
rect 96764 7636 364616 7664
rect 96764 7624 96770 7636
rect 364610 7624 364616 7636
rect 364668 7624 364674 7676
rect 23474 7556 23480 7608
rect 23532 7596 23538 7608
rect 80882 7596 80888 7608
rect 23532 7568 80888 7596
rect 23532 7556 23538 7568
rect 80882 7556 80888 7568
rect 80940 7556 80946 7608
rect 109770 7556 109776 7608
rect 109828 7596 109834 7608
rect 385954 7596 385960 7608
rect 109828 7568 385960 7596
rect 109828 7556 109834 7568
rect 385954 7556 385960 7568
rect 386012 7556 386018 7608
rect 61838 7488 61844 7540
rect 61896 7528 61902 7540
rect 124214 7528 124220 7540
rect 61896 7500 124220 7528
rect 61896 7488 61902 7500
rect 124214 7488 124220 7500
rect 124272 7488 124278 7540
rect 143534 7488 143540 7540
rect 143592 7528 143598 7540
rect 152366 7528 152372 7540
rect 143592 7500 152372 7528
rect 143592 7488 143598 7500
rect 152366 7488 152372 7500
rect 152424 7488 152430 7540
rect 61654 7420 61660 7472
rect 61712 7460 61718 7472
rect 121270 7460 121276 7472
rect 61712 7432 121276 7460
rect 61712 7420 61718 7432
rect 121270 7420 121276 7432
rect 121328 7420 121334 7472
rect 84746 7352 84752 7404
rect 84804 7392 84810 7404
rect 140774 7392 140780 7404
rect 84804 7364 140780 7392
rect 84804 7352 84810 7364
rect 140774 7352 140780 7364
rect 140832 7352 140838 7404
rect 57974 7284 57980 7336
rect 58032 7324 58038 7336
rect 108942 7324 108948 7336
rect 58032 7296 108948 7324
rect 58032 7284 58038 7296
rect 108942 7284 108948 7296
rect 109000 7284 109006 7336
rect 93578 7216 93584 7268
rect 93636 7256 93642 7268
rect 191742 7256 191748 7268
rect 93636 7228 191748 7256
rect 93636 7216 93642 7228
rect 191742 7216 191748 7228
rect 191800 7216 191806 7268
rect 57882 7148 57888 7200
rect 57940 7188 57946 7200
rect 95234 7188 95240 7200
rect 57940 7160 95240 7188
rect 57940 7148 57946 7160
rect 95234 7148 95240 7160
rect 95292 7148 95298 7200
rect 23566 7080 23572 7132
rect 23624 7120 23630 7132
rect 96614 7120 96620 7132
rect 23624 7092 96620 7120
rect 23624 7080 23630 7092
rect 96614 7080 96620 7092
rect 96672 7080 96678 7132
rect 69106 7012 69112 7064
rect 69164 7052 69170 7064
rect 156506 7052 156512 7064
rect 69164 7024 156512 7052
rect 69164 7012 69170 7024
rect 156506 7012 156512 7024
rect 156564 7012 156570 7064
rect 150526 6944 150532 6996
rect 150584 6984 150590 6996
rect 153930 6984 153936 6996
rect 150584 6956 153936 6984
rect 150584 6944 150590 6956
rect 153930 6944 153936 6956
rect 153988 6944 153994 6996
rect 127526 6876 127532 6928
rect 127584 6916 127590 6928
rect 134150 6916 134156 6928
rect 127584 6888 134156 6916
rect 127584 6876 127590 6888
rect 134150 6876 134156 6888
rect 134208 6876 134214 6928
rect 150434 6876 150440 6928
rect 150492 6916 150498 6928
rect 160554 6916 160560 6928
rect 150492 6888 160560 6916
rect 150492 6876 150498 6888
rect 160554 6876 160560 6888
rect 160612 6876 160618 6928
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 17218 6848 17224 6860
rect 3568 6820 17224 6848
rect 3568 6808 3574 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 56594 6808 56600 6860
rect 56652 6848 56658 6860
rect 95418 6848 95424 6860
rect 56652 6820 95424 6848
rect 56652 6808 56658 6820
rect 95418 6808 95424 6820
rect 95476 6808 95482 6860
rect 101398 6808 101404 6860
rect 101456 6848 101462 6860
rect 104894 6848 104900 6860
rect 101456 6820 104900 6848
rect 101456 6808 101462 6820
rect 104894 6808 104900 6820
rect 104952 6808 104958 6860
rect 107562 6808 107568 6860
rect 107620 6848 107626 6860
rect 111150 6848 111156 6860
rect 107620 6820 111156 6848
rect 107620 6808 107626 6820
rect 111150 6808 111156 6820
rect 111208 6808 111214 6860
rect 111518 6808 111524 6860
rect 111576 6848 111582 6860
rect 116026 6848 116032 6860
rect 111576 6820 116032 6848
rect 111576 6808 111582 6820
rect 116026 6808 116032 6820
rect 116084 6808 116090 6860
rect 118694 6808 118700 6860
rect 118752 6848 118758 6860
rect 120994 6848 121000 6860
rect 118752 6820 121000 6848
rect 118752 6808 118758 6820
rect 120994 6808 121000 6820
rect 121052 6808 121058 6860
rect 184750 6808 184756 6860
rect 184808 6848 184814 6860
rect 204806 6848 204812 6860
rect 184808 6820 204812 6848
rect 184808 6808 184814 6820
rect 204806 6808 204812 6820
rect 204864 6808 204870 6860
rect 507210 6808 507216 6860
rect 507268 6848 507274 6860
rect 509602 6848 509608 6860
rect 507268 6820 509608 6848
rect 507268 6808 507274 6820
rect 509602 6808 509608 6820
rect 509660 6808 509666 6860
rect 72878 6740 72884 6792
rect 72936 6780 72942 6792
rect 186314 6780 186320 6792
rect 72936 6752 186320 6780
rect 72936 6740 72942 6752
rect 186314 6740 186320 6752
rect 186372 6740 186378 6792
rect 213730 6740 213736 6792
rect 213788 6780 213794 6792
rect 278682 6780 278688 6792
rect 213788 6752 278688 6780
rect 213788 6740 213794 6752
rect 278682 6740 278688 6752
rect 278740 6740 278746 6792
rect 431402 6740 431408 6792
rect 431460 6780 431466 6792
rect 434622 6780 434628 6792
rect 431460 6752 434628 6780
rect 431460 6740 431466 6752
rect 434622 6740 434628 6752
rect 434680 6740 434686 6792
rect 476022 6740 476028 6792
rect 476080 6780 476086 6792
rect 484854 6780 484860 6792
rect 476080 6752 484860 6780
rect 476080 6740 476086 6752
rect 484854 6740 484860 6752
rect 484912 6740 484918 6792
rect 80882 6672 80888 6724
rect 80940 6712 80946 6724
rect 88334 6712 88340 6724
rect 80940 6684 88340 6712
rect 80940 6672 80946 6684
rect 88334 6672 88340 6684
rect 88392 6672 88398 6724
rect 214558 6712 214564 6724
rect 88444 6684 214564 6712
rect 85114 6604 85120 6656
rect 85172 6644 85178 6656
rect 88444 6644 88472 6684
rect 214558 6672 214564 6684
rect 214616 6672 214622 6724
rect 391842 6672 391848 6724
rect 391900 6712 391906 6724
rect 395430 6712 395436 6724
rect 391900 6684 395436 6712
rect 391900 6672 391906 6684
rect 395430 6672 395436 6684
rect 395488 6672 395494 6724
rect 449158 6672 449164 6724
rect 449216 6712 449222 6724
rect 455690 6712 455696 6724
rect 449216 6684 455696 6712
rect 449216 6672 449222 6684
rect 455690 6672 455696 6684
rect 455748 6672 455754 6724
rect 462314 6672 462320 6724
rect 462372 6712 462378 6724
rect 471054 6712 471060 6724
rect 462372 6684 471060 6712
rect 462372 6672 462378 6684
rect 471054 6672 471060 6684
rect 471112 6672 471118 6724
rect 471974 6672 471980 6724
rect 472032 6712 472038 6724
rect 481726 6712 481732 6724
rect 472032 6684 481732 6712
rect 472032 6672 472038 6684
rect 481726 6672 481732 6684
rect 481784 6672 481790 6724
rect 85172 6616 88472 6644
rect 85172 6604 85178 6616
rect 88610 6604 88616 6656
rect 88668 6644 88674 6656
rect 231762 6644 231768 6656
rect 88668 6616 231768 6644
rect 88668 6604 88674 6616
rect 231762 6604 231768 6616
rect 231820 6604 231826 6656
rect 427722 6604 427728 6656
rect 427780 6644 427786 6656
rect 441522 6644 441528 6656
rect 427780 6616 441528 6644
rect 427780 6604 427786 6616
rect 441522 6604 441528 6616
rect 441580 6604 441586 6656
rect 467098 6604 467104 6656
rect 467156 6644 467162 6656
rect 480530 6644 480536 6656
rect 467156 6616 480536 6644
rect 467156 6604 467162 6616
rect 480530 6604 480536 6616
rect 480588 6604 480594 6656
rect 50614 6536 50620 6588
rect 50672 6576 50678 6588
rect 69106 6576 69112 6588
rect 50672 6548 69112 6576
rect 50672 6536 50678 6548
rect 69106 6536 69112 6548
rect 69164 6536 69170 6588
rect 85574 6536 85580 6588
rect 85632 6576 85638 6588
rect 272518 6576 272524 6588
rect 85632 6548 272524 6576
rect 85632 6536 85638 6548
rect 272518 6536 272524 6548
rect 272576 6536 272582 6588
rect 282822 6536 282828 6588
rect 282880 6576 282886 6588
rect 321554 6576 321560 6588
rect 282880 6548 321560 6576
rect 282880 6536 282886 6548
rect 321554 6536 321560 6548
rect 321612 6536 321618 6588
rect 400122 6536 400128 6588
rect 400180 6576 400186 6588
rect 430850 6576 430856 6588
rect 400180 6548 430856 6576
rect 400180 6536 400186 6548
rect 430850 6536 430856 6548
rect 430908 6536 430914 6588
rect 433978 6536 433984 6588
rect 434036 6576 434042 6588
rect 448514 6576 448520 6588
rect 434036 6548 448520 6576
rect 434036 6536 434042 6548
rect 448514 6536 448520 6548
rect 448572 6536 448578 6588
rect 458082 6536 458088 6588
rect 458140 6576 458146 6588
rect 467558 6576 467564 6588
rect 458140 6548 467564 6576
rect 458140 6536 458146 6548
rect 467558 6536 467564 6548
rect 467616 6536 467622 6588
rect 476758 6536 476764 6588
rect 476816 6576 476822 6588
rect 492306 6576 492312 6588
rect 476816 6548 492312 6576
rect 476816 6536 476822 6548
rect 492306 6536 492312 6548
rect 492364 6536 492370 6588
rect 509878 6536 509884 6588
rect 509936 6576 509942 6588
rect 529014 6576 529020 6588
rect 509936 6548 529020 6576
rect 509936 6536 509942 6548
rect 529014 6536 529020 6548
rect 529072 6536 529078 6588
rect 53098 6468 53104 6520
rect 53156 6508 53162 6520
rect 72602 6508 72608 6520
rect 53156 6480 72608 6508
rect 53156 6468 53162 6480
rect 72602 6468 72608 6480
rect 72660 6468 72666 6520
rect 73890 6468 73896 6520
rect 73948 6508 73954 6520
rect 82078 6508 82084 6520
rect 73948 6480 82084 6508
rect 73948 6468 73954 6480
rect 82078 6468 82084 6480
rect 82136 6468 82142 6520
rect 87230 6468 87236 6520
rect 87288 6508 87294 6520
rect 282914 6508 282920 6520
rect 87288 6480 282920 6508
rect 87288 6468 87294 6480
rect 282914 6468 282920 6480
rect 282972 6468 282978 6520
rect 291746 6468 291752 6520
rect 291804 6508 291810 6520
rect 340138 6508 340144 6520
rect 291804 6480 340144 6508
rect 291804 6468 291810 6480
rect 340138 6468 340144 6480
rect 340196 6468 340202 6520
rect 413094 6508 413100 6520
rect 393286 6480 413100 6508
rect 23014 6400 23020 6452
rect 23072 6440 23078 6452
rect 43070 6440 43076 6452
rect 23072 6412 43076 6440
rect 23072 6400 23078 6412
rect 43070 6400 43076 6412
rect 43128 6400 43134 6452
rect 52270 6400 52276 6452
rect 52328 6440 52334 6452
rect 79686 6440 79692 6452
rect 52328 6412 79692 6440
rect 52328 6400 52334 6412
rect 79686 6400 79692 6412
rect 79744 6400 79750 6452
rect 86310 6400 86316 6452
rect 86368 6440 86374 6452
rect 294966 6440 294972 6452
rect 86368 6412 294972 6440
rect 86368 6400 86374 6412
rect 294966 6400 294972 6412
rect 295024 6400 295030 6452
rect 359550 6400 359556 6452
rect 359608 6440 359614 6452
rect 390646 6440 390652 6452
rect 359608 6412 390652 6440
rect 359608 6400 359614 6412
rect 390646 6400 390652 6412
rect 390704 6400 390710 6452
rect 17678 6332 17684 6384
rect 17736 6372 17742 6384
rect 40310 6372 40316 6384
rect 17736 6344 40316 6372
rect 17736 6332 17742 6344
rect 40310 6332 40316 6344
rect 40368 6332 40374 6384
rect 53374 6332 53380 6384
rect 53432 6372 53438 6384
rect 86862 6372 86868 6384
rect 53432 6344 86868 6372
rect 53432 6332 53438 6344
rect 86862 6332 86868 6344
rect 86920 6332 86926 6384
rect 92198 6332 92204 6384
rect 92256 6372 92262 6384
rect 92256 6344 92520 6372
rect 92256 6332 92262 6344
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 33134 6304 33140 6316
rect 1360 6276 33140 6304
rect 1360 6264 1366 6276
rect 33134 6264 33140 6276
rect 33192 6264 33198 6316
rect 57238 6264 57244 6316
rect 57296 6304 57302 6316
rect 92382 6304 92388 6316
rect 57296 6276 92388 6304
rect 57296 6264 57302 6276
rect 92382 6264 92388 6276
rect 92440 6264 92446 6316
rect 26326 6196 26332 6248
rect 26384 6236 26390 6248
rect 86954 6236 86960 6248
rect 26384 6208 86960 6236
rect 26384 6196 26390 6208
rect 86954 6196 86960 6208
rect 87012 6196 87018 6248
rect 92492 6236 92520 6344
rect 92566 6332 92572 6384
rect 92624 6372 92630 6384
rect 300762 6372 300768 6384
rect 92624 6344 300768 6372
rect 92624 6332 92630 6344
rect 300762 6332 300768 6344
rect 300820 6332 300826 6384
rect 341610 6332 341616 6384
rect 341668 6372 341674 6384
rect 363046 6372 363052 6384
rect 341668 6344 363052 6372
rect 341668 6332 341674 6344
rect 363046 6332 363052 6344
rect 363104 6332 363110 6384
rect 373258 6332 373264 6384
rect 373316 6372 373322 6384
rect 393286 6372 393314 6480
rect 413094 6468 413100 6480
rect 413152 6468 413158 6520
rect 417418 6468 417424 6520
rect 417476 6508 417482 6520
rect 448606 6508 448612 6520
rect 417476 6480 448612 6508
rect 417476 6468 417482 6480
rect 448606 6468 448612 6480
rect 448664 6468 448670 6520
rect 449434 6468 449440 6520
rect 449492 6508 449498 6520
rect 465166 6508 465172 6520
rect 449492 6480 465172 6508
rect 449492 6468 449498 6480
rect 465166 6468 465172 6480
rect 465224 6468 465230 6520
rect 467190 6468 467196 6520
rect 467248 6508 467254 6520
rect 484394 6508 484400 6520
rect 467248 6480 484400 6508
rect 467248 6468 467254 6480
rect 484394 6468 484400 6480
rect 484452 6468 484458 6520
rect 485130 6468 485136 6520
rect 485188 6508 485194 6520
rect 493502 6508 493508 6520
rect 485188 6480 493508 6508
rect 485188 6468 485194 6480
rect 493502 6468 493508 6480
rect 493560 6468 493566 6520
rect 528554 6468 528560 6520
rect 528612 6508 528618 6520
rect 547874 6508 547880 6520
rect 528612 6480 547880 6508
rect 528612 6468 528618 6480
rect 547874 6468 547880 6480
rect 547932 6468 547938 6520
rect 408678 6400 408684 6452
rect 408736 6440 408742 6452
rect 417878 6440 417884 6452
rect 408736 6412 417884 6440
rect 408736 6400 408742 6412
rect 417878 6400 417884 6412
rect 417936 6400 417942 6452
rect 421558 6400 421564 6452
rect 421616 6440 421622 6452
rect 458082 6440 458088 6452
rect 421616 6412 458088 6440
rect 421616 6400 421622 6412
rect 458082 6400 458088 6412
rect 458140 6400 458146 6452
rect 460198 6400 460204 6452
rect 460256 6440 460262 6452
rect 473814 6440 473820 6452
rect 460256 6412 473820 6440
rect 460256 6400 460262 6412
rect 473814 6400 473820 6412
rect 473872 6400 473878 6452
rect 475378 6400 475384 6452
rect 475436 6440 475442 6452
rect 502978 6440 502984 6452
rect 475436 6412 502984 6440
rect 475436 6400 475442 6412
rect 502978 6400 502984 6412
rect 503036 6400 503042 6452
rect 520918 6400 520924 6452
rect 520976 6440 520982 6452
rect 546678 6440 546684 6452
rect 520976 6412 546684 6440
rect 520976 6400 520982 6412
rect 546678 6400 546684 6412
rect 546736 6400 546742 6452
rect 403526 6372 403532 6384
rect 373316 6344 393314 6372
rect 403084 6344 403532 6372
rect 373316 6332 373322 6344
rect 310422 6304 310428 6316
rect 92768 6276 310428 6304
rect 92768 6236 92796 6276
rect 310422 6264 310428 6276
rect 310480 6264 310486 6316
rect 319438 6264 319444 6316
rect 319496 6304 319502 6316
rect 331306 6304 331312 6316
rect 319496 6276 331312 6304
rect 319496 6264 319502 6276
rect 331306 6264 331312 6276
rect 331364 6264 331370 6316
rect 353018 6264 353024 6316
rect 353076 6304 353082 6316
rect 403084 6304 403112 6344
rect 403526 6332 403532 6344
rect 403584 6332 403590 6384
rect 416866 6332 416872 6384
rect 416924 6372 416930 6384
rect 426894 6372 426900 6384
rect 416924 6344 426900 6372
rect 416924 6332 416930 6344
rect 426894 6332 426900 6344
rect 426952 6332 426958 6384
rect 427170 6332 427176 6384
rect 427228 6372 427234 6384
rect 462498 6372 462504 6384
rect 427228 6344 462504 6372
rect 427228 6332 427234 6344
rect 462498 6332 462504 6344
rect 462556 6332 462562 6384
rect 467650 6332 467656 6384
rect 467708 6372 467714 6384
rect 492030 6372 492036 6384
rect 467708 6344 492036 6372
rect 467708 6332 467714 6344
rect 492030 6332 492036 6344
rect 492088 6332 492094 6384
rect 493318 6332 493324 6384
rect 493376 6372 493382 6384
rect 525794 6372 525800 6384
rect 493376 6344 525800 6372
rect 493376 6332 493382 6344
rect 525794 6332 525800 6344
rect 525852 6332 525858 6384
rect 526254 6332 526260 6384
rect 526312 6372 526318 6384
rect 565630 6372 565636 6384
rect 526312 6344 565636 6372
rect 526312 6332 526318 6344
rect 565630 6332 565636 6344
rect 565688 6332 565694 6384
rect 353076 6276 403112 6304
rect 353076 6264 353082 6276
rect 403158 6264 403164 6316
rect 403216 6304 403222 6316
rect 427722 6304 427728 6316
rect 403216 6276 427728 6304
rect 403216 6264 403222 6276
rect 427722 6264 427728 6276
rect 427780 6264 427786 6316
rect 435450 6264 435456 6316
rect 435508 6304 435514 6316
rect 471882 6304 471888 6316
rect 435508 6276 471888 6304
rect 435508 6264 435514 6276
rect 471882 6264 471888 6276
rect 471940 6264 471946 6316
rect 478874 6264 478880 6316
rect 478932 6304 478938 6316
rect 543734 6304 543740 6316
rect 478932 6276 543740 6304
rect 478932 6264 478938 6276
rect 543734 6264 543740 6276
rect 543792 6264 543798 6316
rect 92492 6208 92796 6236
rect 97442 6196 97448 6248
rect 97500 6236 97506 6248
rect 361114 6236 361120 6248
rect 97500 6208 361120 6236
rect 97500 6196 97506 6208
rect 361114 6196 361120 6208
rect 361172 6196 361178 6248
rect 363690 6196 363696 6248
rect 363748 6236 363754 6248
rect 368382 6236 368388 6248
rect 363748 6208 368388 6236
rect 363748 6196 363754 6208
rect 368382 6196 368388 6208
rect 368440 6196 368446 6248
rect 370498 6196 370504 6248
rect 370556 6236 370562 6248
rect 403618 6236 403624 6248
rect 370556 6208 403624 6236
rect 370556 6196 370562 6208
rect 403618 6196 403624 6208
rect 403676 6196 403682 6248
rect 403710 6196 403716 6248
rect 403768 6236 403774 6248
rect 466454 6236 466460 6248
rect 403768 6208 466460 6236
rect 403768 6196 403774 6208
rect 466454 6196 466460 6208
rect 466512 6196 466518 6248
rect 470686 6196 470692 6248
rect 470744 6236 470750 6248
rect 481542 6236 481548 6248
rect 470744 6208 481548 6236
rect 470744 6196 470750 6208
rect 481542 6196 481548 6208
rect 481600 6196 481606 6248
rect 485222 6196 485228 6248
rect 485280 6236 485286 6248
rect 566826 6236 566832 6248
rect 485280 6208 566832 6236
rect 485280 6196 485286 6208
rect 566826 6196 566832 6208
rect 566884 6196 566890 6248
rect 20622 6128 20628 6180
rect 20680 6168 20686 6180
rect 59262 6168 59268 6180
rect 20680 6140 59268 6168
rect 20680 6128 20686 6140
rect 59262 6128 59268 6140
rect 59320 6128 59326 6180
rect 68738 6128 68744 6180
rect 68796 6168 68802 6180
rect 80606 6168 80612 6180
rect 68796 6140 80612 6168
rect 68796 6128 68802 6140
rect 80606 6128 80612 6140
rect 80664 6128 80670 6180
rect 87690 6128 87696 6180
rect 87748 6168 87754 6180
rect 262858 6168 262864 6180
rect 87748 6140 262864 6168
rect 87748 6128 87754 6140
rect 262858 6128 262864 6140
rect 262916 6128 262922 6180
rect 265618 6128 265624 6180
rect 265676 6168 265682 6180
rect 536098 6168 536104 6180
rect 265676 6140 536104 6168
rect 265676 6128 265682 6140
rect 536098 6128 536104 6140
rect 536156 6128 536162 6180
rect 65334 6060 65340 6112
rect 65392 6100 65398 6112
rect 150434 6100 150440 6112
rect 65392 6072 150440 6100
rect 65392 6060 65398 6072
rect 150434 6060 150440 6072
rect 150492 6060 150498 6112
rect 186866 6060 186872 6112
rect 186924 6100 186930 6112
rect 191742 6100 191748 6112
rect 186924 6072 191748 6100
rect 186924 6060 186930 6072
rect 191742 6060 191748 6072
rect 191800 6060 191806 6112
rect 204162 6060 204168 6112
rect 204220 6100 204226 6112
rect 221642 6100 221648 6112
rect 204220 6072 221648 6100
rect 204220 6060 204226 6072
rect 221642 6060 221648 6072
rect 221700 6060 221706 6112
rect 345750 6060 345756 6112
rect 345808 6100 345814 6112
rect 351914 6100 351920 6112
rect 345808 6072 351920 6100
rect 345808 6060 345814 6072
rect 351914 6060 351920 6072
rect 351972 6060 351978 6112
rect 360010 6060 360016 6112
rect 360068 6100 360074 6112
rect 362954 6100 362960 6112
rect 360068 6072 362960 6100
rect 360068 6060 360074 6072
rect 362954 6060 362960 6072
rect 363012 6060 363018 6112
rect 62390 5992 62396 6044
rect 62448 6032 62454 6044
rect 144638 6032 144644 6044
rect 62448 6004 144644 6032
rect 62448 5992 62454 6004
rect 144638 5992 144644 6004
rect 144696 5992 144702 6044
rect 145006 5992 145012 6044
rect 145064 6032 145070 6044
rect 155402 6032 155408 6044
rect 145064 6004 155408 6032
rect 145064 5992 145070 6004
rect 155402 5992 155408 6004
rect 155460 5992 155466 6044
rect 80054 5924 80060 5976
rect 80112 5964 80118 5976
rect 88610 5964 88616 5976
rect 80112 5936 88616 5964
rect 80112 5924 80118 5936
rect 88610 5924 88616 5936
rect 88668 5924 88674 5976
rect 89990 5924 89996 5976
rect 90048 5964 90054 5976
rect 92566 5964 92572 5976
rect 90048 5936 92572 5964
rect 90048 5924 90054 5936
rect 92566 5924 92572 5936
rect 92624 5924 92630 5976
rect 127618 5924 127624 5976
rect 127676 5964 127682 5976
rect 140682 5964 140688 5976
rect 127676 5936 140688 5964
rect 127676 5924 127682 5936
rect 140682 5924 140688 5936
rect 140740 5924 140746 5976
rect 94498 5856 94504 5908
rect 94556 5896 94562 5908
rect 97994 5896 98000 5908
rect 94556 5868 98000 5896
rect 94556 5856 94562 5868
rect 97994 5856 98000 5868
rect 98052 5856 98058 5908
rect 140130 5856 140136 5908
rect 140188 5896 140194 5908
rect 146662 5896 146668 5908
rect 140188 5868 146668 5896
rect 140188 5856 140194 5868
rect 146662 5856 146668 5868
rect 146720 5856 146726 5908
rect 66990 5788 66996 5840
rect 67048 5828 67054 5840
rect 174262 5828 174268 5840
rect 67048 5800 174268 5828
rect 67048 5788 67054 5800
rect 174262 5788 174268 5800
rect 174320 5788 174326 5840
rect 367830 5652 367836 5704
rect 367888 5692 367894 5704
rect 370958 5692 370964 5704
rect 367888 5664 370964 5692
rect 367888 5652 367894 5664
rect 370958 5652 370964 5664
rect 371016 5652 371022 5704
rect 151078 5624 151084 5636
rect 149072 5596 151084 5624
rect 59630 5516 59636 5568
rect 59688 5556 59694 5568
rect 67542 5556 67548 5568
rect 59688 5528 67548 5556
rect 59688 5516 59694 5528
rect 67542 5516 67548 5528
rect 67600 5516 67606 5568
rect 83182 5448 83188 5500
rect 83240 5488 83246 5500
rect 86678 5488 86684 5500
rect 83240 5460 86684 5488
rect 83240 5448 83246 5460
rect 86678 5448 86684 5460
rect 86736 5448 86742 5500
rect 86954 5448 86960 5500
rect 87012 5488 87018 5500
rect 97350 5488 97356 5500
rect 87012 5460 97356 5488
rect 87012 5448 87018 5460
rect 97350 5448 97356 5460
rect 97408 5448 97414 5500
rect 103514 5448 103520 5500
rect 103572 5488 103578 5500
rect 109218 5488 109224 5500
rect 103572 5460 109224 5488
rect 103572 5448 103578 5460
rect 109218 5448 109224 5460
rect 109276 5448 109282 5500
rect 113266 5448 113272 5500
rect 113324 5488 113330 5500
rect 116394 5488 116400 5500
rect 113324 5460 116400 5488
rect 113324 5448 113330 5460
rect 116394 5448 116400 5460
rect 116452 5448 116458 5500
rect 144730 5448 144736 5500
rect 144788 5488 144794 5500
rect 149072 5488 149100 5596
rect 151078 5584 151084 5596
rect 151136 5584 151142 5636
rect 454770 5584 454776 5636
rect 454828 5624 454834 5636
rect 459554 5624 459560 5636
rect 454828 5596 459560 5624
rect 454828 5584 454834 5596
rect 459554 5584 459560 5596
rect 459612 5584 459618 5636
rect 150434 5516 150440 5568
rect 150492 5556 150498 5568
rect 154298 5556 154304 5568
rect 150492 5528 154304 5556
rect 150492 5516 150498 5528
rect 154298 5516 154304 5528
rect 154356 5516 154362 5568
rect 277394 5516 277400 5568
rect 277452 5556 277458 5568
rect 283098 5556 283104 5568
rect 277452 5528 283104 5556
rect 277452 5516 277458 5528
rect 283098 5516 283104 5528
rect 283156 5516 283162 5568
rect 314010 5516 314016 5568
rect 314068 5556 314074 5568
rect 316218 5556 316224 5568
rect 314068 5528 316224 5556
rect 314068 5516 314074 5528
rect 316218 5516 316224 5528
rect 316276 5516 316282 5568
rect 394694 5516 394700 5568
rect 394752 5556 394758 5568
rect 400122 5556 400128 5568
rect 394752 5528 400128 5556
rect 394752 5516 394758 5528
rect 400122 5516 400128 5528
rect 400180 5516 400186 5568
rect 412634 5516 412640 5568
rect 412692 5556 412698 5568
rect 415486 5556 415492 5568
rect 412692 5528 415492 5556
rect 412692 5516 412698 5528
rect 415486 5516 415492 5528
rect 415544 5516 415550 5568
rect 454678 5516 454684 5568
rect 454736 5556 454742 5568
rect 462774 5556 462780 5568
rect 454736 5528 462780 5556
rect 454736 5516 454742 5528
rect 462774 5516 462780 5528
rect 462832 5516 462838 5568
rect 471238 5516 471244 5568
rect 471296 5556 471302 5568
rect 476942 5556 476948 5568
rect 471296 5528 476948 5556
rect 471296 5516 471302 5528
rect 476942 5516 476948 5528
rect 477000 5516 477006 5568
rect 491294 5516 491300 5568
rect 491352 5556 491358 5568
rect 494698 5556 494704 5568
rect 491352 5528 494704 5556
rect 491352 5516 491358 5528
rect 494698 5516 494704 5528
rect 494756 5516 494762 5568
rect 534810 5516 534816 5568
rect 534868 5556 534874 5568
rect 539594 5556 539600 5568
rect 534868 5528 539600 5556
rect 534868 5516 534874 5528
rect 539594 5516 539600 5528
rect 539652 5516 539658 5568
rect 144788 5460 149100 5488
rect 144788 5448 144794 5460
rect 149146 5448 149152 5500
rect 149204 5488 149210 5500
rect 155218 5488 155224 5500
rect 149204 5460 155224 5488
rect 149204 5448 149210 5460
rect 155218 5448 155224 5460
rect 155276 5448 155282 5500
rect 180150 5448 180156 5500
rect 180208 5488 180214 5500
rect 185026 5488 185032 5500
rect 180208 5460 185032 5488
rect 180208 5448 180214 5460
rect 185026 5448 185032 5460
rect 185084 5448 185090 5500
rect 84378 5380 84384 5432
rect 84436 5420 84442 5432
rect 179414 5420 179420 5432
rect 84436 5392 179420 5420
rect 84436 5380 84442 5392
rect 179414 5380 179420 5392
rect 179472 5380 179478 5432
rect 71958 5312 71964 5364
rect 72016 5352 72022 5364
rect 198826 5352 198832 5364
rect 72016 5324 198832 5352
rect 72016 5312 72022 5324
rect 198826 5312 198832 5324
rect 198884 5312 198890 5364
rect 232038 5312 232044 5364
rect 232096 5352 232102 5364
rect 247586 5352 247592 5364
rect 232096 5324 247592 5352
rect 232096 5312 232102 5324
rect 247586 5312 247592 5324
rect 247644 5312 247650 5364
rect 59446 5244 59452 5296
rect 59504 5284 59510 5296
rect 60918 5284 60924 5296
rect 59504 5256 60924 5284
rect 59504 5244 59510 5256
rect 60918 5244 60924 5256
rect 60976 5244 60982 5296
rect 79410 5244 79416 5296
rect 79468 5284 79474 5296
rect 212994 5284 213000 5296
rect 79468 5256 213000 5284
rect 79468 5244 79474 5256
rect 212994 5244 213000 5256
rect 213052 5244 213058 5296
rect 214558 5244 214564 5296
rect 214616 5284 214622 5296
rect 235994 5284 236000 5296
rect 214616 5256 236000 5284
rect 214616 5244 214622 5256
rect 235994 5244 236000 5256
rect 236052 5244 236058 5296
rect 74166 5176 74172 5228
rect 74224 5216 74230 5228
rect 205634 5216 205640 5228
rect 74224 5188 205640 5216
rect 74224 5176 74230 5188
rect 205634 5176 205640 5188
rect 205692 5176 205698 5228
rect 207658 5176 207664 5228
rect 207716 5216 207722 5228
rect 346946 5216 346952 5228
rect 207716 5188 346952 5216
rect 207716 5176 207722 5188
rect 346946 5176 346952 5188
rect 347004 5176 347010 5228
rect 51810 5108 51816 5160
rect 51868 5148 51874 5160
rect 66714 5148 66720 5160
rect 51868 5120 66720 5148
rect 51868 5108 51874 5120
rect 66714 5108 66720 5120
rect 66772 5108 66778 5160
rect 82998 5108 83004 5160
rect 83056 5148 83062 5160
rect 224954 5148 224960 5160
rect 83056 5120 224960 5148
rect 83056 5108 83062 5120
rect 224954 5108 224960 5120
rect 225012 5108 225018 5160
rect 236362 5108 236368 5160
rect 236420 5148 236426 5160
rect 315022 5148 315028 5160
rect 236420 5120 315028 5148
rect 236420 5108 236426 5120
rect 315022 5108 315028 5120
rect 315080 5108 315086 5160
rect 55858 5040 55864 5092
rect 55916 5080 55922 5092
rect 80882 5080 80888 5092
rect 55916 5052 80888 5080
rect 55916 5040 55922 5052
rect 80882 5040 80888 5052
rect 80940 5040 80946 5092
rect 84654 5040 84660 5092
rect 84712 5080 84718 5092
rect 274634 5080 274640 5092
rect 84712 5052 274640 5080
rect 84712 5040 84718 5052
rect 274634 5040 274640 5052
rect 274692 5040 274698 5092
rect 51902 4972 51908 5024
rect 51960 5012 51966 5024
rect 77386 5012 77392 5024
rect 51960 4984 77392 5012
rect 51960 4972 51966 4984
rect 77386 4972 77392 4984
rect 77444 4972 77450 5024
rect 88518 4972 88524 5024
rect 88576 5012 88582 5024
rect 291746 5012 291752 5024
rect 88576 4984 291752 5012
rect 88576 4972 88582 4984
rect 291746 4972 291752 4984
rect 291804 4972 291810 5024
rect 27706 4904 27712 4956
rect 27764 4944 27770 4956
rect 44358 4944 44364 4956
rect 27764 4916 44364 4944
rect 27764 4904 27770 4916
rect 44358 4904 44364 4916
rect 44416 4904 44422 4956
rect 53006 4904 53012 4956
rect 53064 4944 53070 4956
rect 84470 4944 84476 4956
rect 53064 4916 84476 4944
rect 53064 4904 53070 4916
rect 84470 4904 84476 4916
rect 84528 4904 84534 4956
rect 86770 4904 86776 4956
rect 86828 4944 86834 4956
rect 301958 4944 301964 4956
rect 86828 4916 301964 4944
rect 86828 4904 86834 4916
rect 301958 4904 301964 4916
rect 302016 4904 302022 4956
rect 11146 4836 11152 4888
rect 11204 4876 11210 4888
rect 41690 4876 41696 4888
rect 11204 4848 41696 4876
rect 11204 4836 11210 4848
rect 41690 4836 41696 4848
rect 41748 4836 41754 4888
rect 54938 4836 54944 4888
rect 54996 4876 55002 4888
rect 87966 4876 87972 4888
rect 54996 4848 87972 4876
rect 54996 4836 55002 4848
rect 87966 4836 87972 4848
rect 88024 4836 88030 4888
rect 109678 4836 109684 4888
rect 109736 4876 109742 4888
rect 111794 4876 111800 4888
rect 109736 4848 111800 4876
rect 109736 4836 109742 4848
rect 111794 4836 111800 4848
rect 111852 4836 111858 4888
rect 114462 4836 114468 4888
rect 114520 4876 114526 4888
rect 118050 4876 118056 4888
rect 114520 4848 118056 4876
rect 114520 4836 114526 4848
rect 118050 4836 118056 4848
rect 118108 4836 118114 4888
rect 121178 4836 121184 4888
rect 121236 4876 121242 4888
rect 489914 4876 489920 4888
rect 121236 4848 489920 4876
rect 121236 4836 121242 4848
rect 489914 4836 489920 4848
rect 489972 4836 489978 4888
rect 22738 4768 22744 4820
rect 22796 4808 22802 4820
rect 56502 4808 56508 4820
rect 22796 4780 56508 4808
rect 22796 4768 22802 4780
rect 56502 4768 56508 4780
rect 56560 4768 56566 4820
rect 68554 4768 68560 4820
rect 68612 4808 68618 4820
rect 68612 4780 74534 4808
rect 68612 4768 68618 4780
rect 56042 4700 56048 4752
rect 56100 4740 56106 4752
rect 73798 4740 73804 4752
rect 56100 4712 73804 4740
rect 56100 4700 56106 4712
rect 73798 4700 73804 4712
rect 73856 4700 73862 4752
rect 74506 4740 74534 4780
rect 108390 4768 108396 4820
rect 108448 4808 108454 4820
rect 114094 4808 114100 4820
rect 108448 4780 114100 4808
rect 108448 4768 108454 4780
rect 114094 4768 114100 4780
rect 114152 4768 114158 4820
rect 121454 4768 121460 4820
rect 121512 4808 121518 4820
rect 521562 4808 521568 4820
rect 121512 4780 521568 4808
rect 121512 4768 121518 4780
rect 521562 4768 521568 4780
rect 521620 4768 521626 4820
rect 139394 4740 139400 4752
rect 74506 4712 139400 4740
rect 139394 4700 139400 4712
rect 139452 4700 139458 4752
rect 146570 4700 146576 4752
rect 146628 4740 146634 4752
rect 149146 4740 149152 4752
rect 146628 4712 149152 4740
rect 146628 4700 146634 4712
rect 149146 4700 149152 4712
rect 149204 4700 149210 4752
rect 68646 4632 68652 4684
rect 68704 4672 68710 4684
rect 133782 4672 133788 4684
rect 68704 4644 133788 4672
rect 68704 4632 68710 4644
rect 133782 4632 133788 4644
rect 133840 4632 133846 4684
rect 76190 4564 76196 4616
rect 76248 4604 76254 4616
rect 127618 4604 127624 4616
rect 76248 4576 127624 4604
rect 76248 4564 76254 4576
rect 127618 4564 127624 4576
rect 127676 4564 127682 4616
rect 131114 4564 131120 4616
rect 131172 4604 131178 4616
rect 137922 4604 137928 4616
rect 131172 4576 137928 4604
rect 131172 4564 131178 4576
rect 137922 4564 137928 4576
rect 137980 4564 137986 4616
rect 59262 4496 59268 4548
rect 59320 4536 59326 4548
rect 101674 4536 101680 4548
rect 59320 4508 101680 4536
rect 59320 4496 59326 4508
rect 101674 4496 101680 4508
rect 101732 4496 101738 4548
rect 62574 4428 62580 4480
rect 62632 4468 62638 4480
rect 62632 4440 142154 4468
rect 62632 4428 62638 4440
rect 142126 4196 142154 4440
rect 153746 4360 153752 4412
rect 153804 4400 153810 4412
rect 156598 4400 156604 4412
rect 153804 4372 156604 4400
rect 153804 4360 153810 4372
rect 156598 4360 156604 4372
rect 156656 4360 156662 4412
rect 144822 4224 144828 4276
rect 144880 4264 144886 4276
rect 150526 4264 150532 4276
rect 144880 4236 150532 4264
rect 144880 4224 144886 4236
rect 150526 4224 150532 4236
rect 150584 4224 150590 4276
rect 142126 4168 144868 4196
rect 54570 4088 54576 4140
rect 54628 4128 54634 4140
rect 57238 4128 57244 4140
rect 54628 4100 57244 4128
rect 54628 4088 54634 4100
rect 57238 4088 57244 4100
rect 57296 4088 57302 4140
rect 75178 4088 75184 4140
rect 75236 4128 75242 4140
rect 106918 4128 106924 4140
rect 75236 4100 106924 4128
rect 75236 4088 75242 4100
rect 106918 4088 106924 4100
rect 106976 4088 106982 4140
rect 109494 4088 109500 4140
rect 109552 4128 109558 4140
rect 116670 4128 116676 4140
rect 109552 4100 116676 4128
rect 109552 4088 109558 4100
rect 116670 4088 116676 4100
rect 116728 4088 116734 4140
rect 119430 4088 119436 4140
rect 119488 4128 119494 4140
rect 123478 4128 123484 4140
rect 119488 4100 123484 4128
rect 119488 4088 119494 4100
rect 123478 4088 123484 4100
rect 123536 4088 123542 4140
rect 127618 4088 127624 4140
rect 127676 4128 127682 4140
rect 131114 4128 131120 4140
rect 127676 4100 131120 4128
rect 127676 4088 127682 4100
rect 131114 4088 131120 4100
rect 131172 4088 131178 4140
rect 144840 4128 144868 4168
rect 145926 4128 145932 4140
rect 144840 4100 145932 4128
rect 145926 4088 145932 4100
rect 145984 4088 145990 4140
rect 251818 4088 251824 4140
rect 251876 4128 251882 4140
rect 252462 4128 252468 4140
rect 251876 4100 252468 4128
rect 251876 4088 251882 4100
rect 252462 4088 252468 4100
rect 252520 4088 252526 4140
rect 313918 4088 313924 4140
rect 313976 4128 313982 4140
rect 317322 4128 317328 4140
rect 313976 4100 317328 4128
rect 313976 4088 313982 4100
rect 317322 4088 317328 4100
rect 317380 4088 317386 4140
rect 362954 4088 362960 4140
rect 363012 4128 363018 4140
rect 367002 4128 367008 4140
rect 363012 4100 367008 4128
rect 363012 4088 363018 4100
rect 367002 4088 367008 4100
rect 367060 4088 367066 4140
rect 516778 4088 516784 4140
rect 516836 4128 516842 4140
rect 519538 4128 519544 4140
rect 516836 4100 519544 4128
rect 516836 4088 516842 4100
rect 519538 4088 519544 4100
rect 519596 4088 519602 4140
rect 59170 4020 59176 4072
rect 59228 4060 59234 4072
rect 124674 4060 124680 4072
rect 59228 4032 124680 4060
rect 59228 4020 59234 4032
rect 124674 4020 124680 4032
rect 124732 4020 124738 4072
rect 127802 4020 127808 4072
rect 127860 4060 127866 4072
rect 137646 4060 137652 4072
rect 127860 4032 137652 4060
rect 127860 4020 127866 4032
rect 137646 4020 137652 4032
rect 137704 4020 137710 4072
rect 146938 4020 146944 4072
rect 146996 4060 147002 4072
rect 157978 4060 157984 4072
rect 146996 4032 157984 4060
rect 146996 4020 147002 4032
rect 157978 4020 157984 4032
rect 158036 4020 158042 4072
rect 180058 4020 180064 4072
rect 180116 4060 180122 4072
rect 187326 4060 187332 4072
rect 180116 4032 187332 4060
rect 180116 4020 180122 4032
rect 187326 4020 187332 4032
rect 187384 4020 187390 4072
rect 85022 3952 85028 4004
rect 85080 3992 85086 4004
rect 156598 3992 156604 4004
rect 85080 3964 156604 3992
rect 85080 3952 85086 3964
rect 156598 3952 156604 3964
rect 156656 3952 156662 4004
rect 179414 3952 179420 4004
rect 179472 3992 179478 4004
rect 192018 3992 192024 4004
rect 179472 3964 192024 3992
rect 179472 3952 179478 3964
rect 192018 3952 192024 3964
rect 192076 3952 192082 4004
rect 234522 3952 234528 4004
rect 234580 3992 234586 4004
rect 251174 3992 251180 4004
rect 234580 3964 251180 3992
rect 234580 3952 234586 3964
rect 251174 3952 251180 3964
rect 251232 3952 251238 4004
rect 460290 3952 460296 4004
rect 460348 3992 460354 4004
rect 469858 3992 469864 4004
rect 460348 3964 469864 3992
rect 460348 3952 460354 3964
rect 469858 3952 469864 3964
rect 469916 3952 469922 4004
rect 71130 3884 71136 3936
rect 71188 3924 71194 3936
rect 152918 3924 152924 3936
rect 71188 3896 152924 3924
rect 71188 3884 71194 3896
rect 152918 3884 152924 3896
rect 152976 3884 152982 3936
rect 172514 3884 172520 3936
rect 172572 3924 172578 3936
rect 181438 3924 181444 3936
rect 172572 3896 181444 3924
rect 172572 3884 172578 3896
rect 181438 3884 181444 3896
rect 181496 3884 181502 3936
rect 186314 3884 186320 3936
rect 186372 3924 186378 3936
rect 212166 3924 212172 3936
rect 186372 3896 212172 3924
rect 186372 3884 186378 3896
rect 212166 3884 212172 3896
rect 212224 3884 212230 3936
rect 212994 3884 213000 3936
rect 213052 3924 213058 3936
rect 238110 3924 238116 3936
rect 213052 3896 238116 3924
rect 213052 3884 213058 3896
rect 238110 3884 238116 3896
rect 238168 3884 238174 3936
rect 240778 3884 240784 3936
rect 240836 3924 240842 3936
rect 244182 3924 244188 3936
rect 240836 3896 244188 3924
rect 240836 3884 240842 3896
rect 244182 3884 244188 3896
rect 244240 3884 244246 3936
rect 262858 3884 262864 3936
rect 262916 3924 262922 3936
rect 262916 3896 267734 3924
rect 262916 3884 262922 3896
rect 33594 3816 33600 3868
rect 33652 3856 33658 3868
rect 36538 3856 36544 3868
rect 33652 3828 36544 3856
rect 33652 3816 33658 3828
rect 36538 3816 36544 3828
rect 36596 3816 36602 3868
rect 43070 3816 43076 3868
rect 43128 3856 43134 3868
rect 46566 3856 46572 3868
rect 43128 3828 46572 3856
rect 43128 3816 43134 3828
rect 46566 3816 46572 3828
rect 46624 3816 46630 3868
rect 61562 3816 61568 3868
rect 61620 3856 61626 3868
rect 85666 3856 85672 3868
rect 61620 3828 85672 3856
rect 61620 3816 61626 3828
rect 85666 3816 85672 3828
rect 85724 3816 85730 3868
rect 90174 3816 90180 3868
rect 90232 3856 90238 3868
rect 92750 3856 92756 3868
rect 90232 3828 92756 3856
rect 90232 3816 90238 3828
rect 92750 3816 92756 3828
rect 92808 3816 92814 3868
rect 93854 3816 93860 3868
rect 93912 3856 93918 3868
rect 97442 3856 97448 3868
rect 93912 3828 97448 3856
rect 93912 3816 93918 3828
rect 97442 3816 97448 3828
rect 97500 3816 97506 3868
rect 101214 3816 101220 3868
rect 101272 3856 101278 3868
rect 101272 3828 103468 3856
rect 101272 3816 101278 3828
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 45278 3788 45284 3800
rect 34848 3760 45284 3788
rect 34848 3748 34854 3760
rect 45278 3748 45284 3760
rect 45336 3748 45342 3800
rect 49510 3748 49516 3800
rect 49568 3788 49574 3800
rect 62022 3788 62028 3800
rect 49568 3760 62028 3788
rect 49568 3748 49574 3760
rect 62022 3748 62028 3760
rect 62080 3748 62086 3800
rect 64138 3748 64144 3800
rect 64196 3788 64202 3800
rect 69658 3788 69664 3800
rect 64196 3760 69664 3788
rect 64196 3748 64202 3760
rect 69658 3748 69664 3760
rect 69716 3748 69722 3800
rect 73890 3748 73896 3800
rect 73948 3788 73954 3800
rect 101030 3788 101036 3800
rect 73948 3760 101036 3788
rect 73948 3748 73954 3760
rect 101030 3748 101036 3760
rect 101088 3748 101094 3800
rect 103440 3788 103468 3828
rect 104250 3816 104256 3868
rect 104308 3856 104314 3868
rect 108390 3856 108396 3868
rect 104308 3828 108396 3856
rect 104308 3816 104314 3828
rect 108390 3816 108396 3828
rect 108448 3816 108454 3868
rect 108574 3816 108580 3868
rect 108632 3856 108638 3868
rect 195974 3856 195980 3868
rect 108632 3828 195980 3856
rect 108632 3816 108638 3828
rect 195974 3816 195980 3828
rect 196032 3816 196038 3868
rect 198826 3816 198832 3868
rect 198884 3856 198890 3868
rect 198884 3828 205588 3856
rect 198884 3816 198890 3828
rect 108206 3788 108212 3800
rect 103440 3760 108212 3788
rect 108206 3748 108212 3760
rect 108264 3748 108270 3800
rect 108482 3748 108488 3800
rect 108540 3788 108546 3800
rect 201678 3788 201684 3800
rect 108540 3760 201684 3788
rect 108540 3748 108546 3760
rect 201678 3748 201684 3760
rect 201736 3748 201742 3800
rect 205560 3788 205588 3828
rect 205634 3816 205640 3868
rect 205692 3856 205698 3868
rect 220446 3856 220452 3868
rect 205692 3828 220452 3856
rect 205692 3816 205698 3828
rect 220446 3816 220452 3828
rect 220504 3816 220510 3868
rect 231762 3816 231768 3868
rect 231820 3856 231826 3868
rect 258258 3856 258264 3868
rect 231820 3828 258264 3856
rect 231820 3816 231826 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 261478 3816 261484 3868
rect 261536 3856 261542 3868
rect 266538 3856 266544 3868
rect 261536 3828 266544 3856
rect 261536 3816 261542 3828
rect 266538 3816 266544 3828
rect 266596 3816 266602 3868
rect 267706 3856 267734 3896
rect 278682 3884 278688 3936
rect 278740 3924 278746 3936
rect 278740 3896 287054 3924
rect 278740 3884 278746 3896
rect 273622 3856 273628 3868
rect 267706 3828 273628 3856
rect 273622 3816 273628 3828
rect 273680 3816 273686 3868
rect 282914 3816 282920 3868
rect 282972 3856 282978 3868
rect 285122 3856 285128 3868
rect 282972 3828 285128 3856
rect 282972 3816 282978 3828
rect 285122 3816 285128 3828
rect 285180 3816 285186 3868
rect 287026 3856 287054 3896
rect 305638 3884 305644 3936
rect 305696 3924 305702 3936
rect 313826 3924 313832 3936
rect 305696 3896 313832 3924
rect 305696 3884 305702 3896
rect 313826 3884 313832 3896
rect 313884 3884 313890 3936
rect 459554 3884 459560 3936
rect 459612 3924 459618 3936
rect 467466 3924 467472 3936
rect 459612 3896 467472 3924
rect 459612 3884 459618 3896
rect 467466 3884 467472 3896
rect 467524 3884 467530 3936
rect 467558 3884 467564 3936
rect 467616 3924 467622 3936
rect 479334 3924 479340 3936
rect 467616 3896 479340 3924
rect 467616 3884 467622 3896
rect 479334 3884 479340 3896
rect 479392 3884 479398 3936
rect 291378 3856 291384 3868
rect 287026 3828 291384 3856
rect 291378 3816 291384 3828
rect 291436 3816 291442 3868
rect 292206 3816 292212 3868
rect 292264 3856 292270 3868
rect 307938 3856 307944 3868
rect 292264 3828 307944 3856
rect 292264 3816 292270 3828
rect 307938 3816 307944 3828
rect 307996 3816 308002 3868
rect 309870 3816 309876 3868
rect 309928 3856 309934 3868
rect 325602 3856 325608 3868
rect 309928 3828 325608 3856
rect 309928 3816 309934 3828
rect 325602 3816 325608 3828
rect 325660 3816 325666 3868
rect 330846 3816 330852 3868
rect 330904 3856 330910 3868
rect 339862 3856 339868 3868
rect 330904 3828 339868 3856
rect 330904 3816 330910 3828
rect 339862 3816 339868 3828
rect 339920 3816 339926 3868
rect 342070 3816 342076 3868
rect 342128 3856 342134 3868
rect 348050 3856 348056 3868
rect 342128 3828 348056 3856
rect 342128 3816 342134 3828
rect 348050 3816 348056 3828
rect 348108 3816 348114 3868
rect 448514 3816 448520 3868
rect 448572 3856 448578 3868
rect 474550 3856 474556 3868
rect 448572 3828 474556 3856
rect 448572 3816 448578 3828
rect 474550 3816 474556 3828
rect 474608 3816 474614 3868
rect 494790 3816 494796 3868
rect 494848 3856 494854 3868
rect 507670 3856 507676 3868
rect 494848 3828 507676 3856
rect 494848 3816 494854 3828
rect 507670 3816 507676 3828
rect 507728 3816 507734 3868
rect 206186 3788 206192 3800
rect 205560 3760 206192 3788
rect 206186 3748 206192 3760
rect 206244 3748 206250 3800
rect 211798 3748 211804 3800
rect 211856 3788 211862 3800
rect 227530 3788 227536 3800
rect 211856 3760 227536 3788
rect 211856 3748 211862 3760
rect 227530 3748 227536 3760
rect 227588 3748 227594 3800
rect 235994 3748 236000 3800
rect 236052 3788 236058 3800
rect 276106 3788 276112 3800
rect 236052 3760 276112 3788
rect 236052 3748 236058 3760
rect 276106 3748 276112 3760
rect 276164 3748 276170 3800
rect 276658 3748 276664 3800
rect 276716 3788 276722 3800
rect 290182 3788 290188 3800
rect 276716 3760 290188 3788
rect 276716 3748 276722 3760
rect 290182 3748 290188 3760
rect 290240 3748 290246 3800
rect 291746 3748 291752 3800
rect 291804 3788 291810 3800
rect 311434 3788 311440 3800
rect 291804 3760 311440 3788
rect 291804 3748 291810 3760
rect 311434 3748 311440 3760
rect 311492 3748 311498 3800
rect 321554 3748 321560 3800
rect 321612 3788 321618 3800
rect 321612 3760 331260 3788
rect 321612 3748 321618 3760
rect 43438 3720 43444 3732
rect 39684 3692 43444 3720
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 39684 3584 39712 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 48958 3680 48964 3732
rect 49016 3720 49022 3732
rect 49016 3692 55214 3720
rect 49016 3680 49022 3692
rect 40678 3612 40684 3664
rect 40736 3652 40742 3664
rect 40736 3624 45554 3652
rect 40736 3612 40742 3624
rect 32456 3556 39712 3584
rect 32456 3544 32462 3556
rect 41874 3544 41880 3596
rect 41932 3584 41938 3596
rect 44818 3584 44824 3596
rect 41932 3556 44824 3584
rect 41932 3544 41938 3556
rect 44818 3544 44824 3556
rect 44876 3544 44882 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 13078 3516 13084 3528
rect 12400 3488 13084 3516
rect 12400 3476 12406 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 42150 3516 42156 3528
rect 38436 3488 42156 3516
rect 38436 3476 38442 3488
rect 42150 3476 42156 3488
rect 42208 3476 42214 3528
rect 45526 3516 45554 3624
rect 49326 3612 49332 3664
rect 49384 3652 49390 3664
rect 55186 3652 55214 3692
rect 57330 3680 57336 3732
rect 57388 3720 57394 3732
rect 89162 3720 89168 3732
rect 57388 3692 89168 3720
rect 57388 3680 57394 3692
rect 89162 3680 89168 3692
rect 89220 3680 89226 3732
rect 92474 3680 92480 3732
rect 92532 3720 92538 3732
rect 93946 3720 93952 3732
rect 92532 3692 93952 3720
rect 92532 3680 92538 3692
rect 93946 3680 93952 3692
rect 94004 3680 94010 3732
rect 103330 3720 103336 3732
rect 94424 3692 103336 3720
rect 58434 3652 58440 3664
rect 49384 3624 52684 3652
rect 55186 3624 58440 3652
rect 49384 3612 49390 3624
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 52546 3584 52552 3596
rect 50580 3556 52552 3584
rect 50580 3544 50586 3556
rect 52546 3544 52552 3556
rect 52604 3544 52610 3596
rect 52656 3584 52684 3624
rect 58434 3612 58440 3624
rect 58492 3612 58498 3664
rect 61378 3612 61384 3664
rect 61436 3652 61442 3664
rect 92934 3652 92940 3664
rect 61436 3624 92940 3652
rect 61436 3612 61442 3624
rect 92934 3612 92940 3624
rect 92992 3612 92998 3664
rect 60826 3584 60832 3596
rect 52656 3556 60832 3584
rect 60826 3544 60832 3556
rect 60884 3544 60890 3596
rect 66898 3544 66904 3596
rect 66956 3584 66962 3596
rect 94424 3584 94452 3692
rect 103330 3680 103336 3692
rect 103388 3680 103394 3732
rect 103422 3680 103428 3732
rect 103480 3720 103486 3732
rect 200666 3720 200672 3732
rect 103480 3692 200672 3720
rect 103480 3680 103486 3692
rect 200666 3680 200672 3692
rect 200724 3680 200730 3732
rect 204806 3680 204812 3732
rect 204864 3720 204870 3732
rect 233418 3720 233424 3732
rect 204864 3692 233424 3720
rect 204864 3680 204870 3692
rect 233418 3680 233424 3692
rect 233476 3680 233482 3732
rect 242894 3680 242900 3732
rect 242952 3720 242958 3732
rect 244090 3720 244096 3732
rect 242952 3692 244096 3720
rect 242952 3680 242958 3692
rect 244090 3680 244096 3692
rect 244148 3680 244154 3732
rect 244182 3680 244188 3732
rect 244240 3720 244246 3732
rect 248782 3720 248788 3732
rect 244240 3692 248788 3720
rect 244240 3680 244246 3692
rect 248782 3680 248788 3692
rect 248840 3680 248846 3732
rect 249058 3680 249064 3732
rect 249116 3720 249122 3732
rect 272426 3720 272432 3732
rect 249116 3692 272432 3720
rect 249116 3680 249122 3692
rect 272426 3680 272432 3692
rect 272484 3680 272490 3732
rect 272518 3680 272524 3732
rect 272576 3720 272582 3732
rect 293678 3720 293684 3732
rect 272576 3692 293684 3720
rect 272576 3680 272582 3692
rect 293678 3680 293684 3692
rect 293736 3680 293742 3732
rect 300762 3680 300768 3732
rect 300820 3720 300826 3732
rect 322106 3720 322112 3732
rect 300820 3692 322112 3720
rect 300820 3680 300826 3692
rect 322106 3680 322112 3692
rect 322164 3680 322170 3732
rect 327718 3680 327724 3732
rect 327776 3720 327782 3732
rect 330386 3720 330392 3732
rect 327776 3692 330392 3720
rect 327776 3680 327782 3692
rect 330386 3680 330392 3692
rect 330444 3680 330450 3732
rect 331232 3720 331260 3760
rect 331306 3748 331312 3800
rect 331364 3788 331370 3800
rect 342162 3788 342168 3800
rect 331364 3760 342168 3788
rect 331364 3748 331370 3760
rect 342162 3748 342168 3760
rect 342220 3748 342226 3800
rect 452654 3748 452660 3800
rect 452712 3788 452718 3800
rect 466270 3788 466276 3800
rect 452712 3760 466276 3788
rect 452712 3748 452718 3760
rect 466270 3748 466276 3760
rect 466328 3748 466334 3800
rect 466454 3748 466460 3800
rect 466512 3788 466518 3800
rect 497090 3788 497096 3800
rect 466512 3760 497096 3788
rect 466512 3748 466518 3760
rect 497090 3748 497096 3760
rect 497148 3748 497154 3800
rect 333882 3720 333888 3732
rect 331232 3692 333888 3720
rect 333882 3680 333888 3692
rect 333940 3680 333946 3732
rect 334618 3680 334624 3732
rect 334676 3720 334682 3732
rect 344554 3720 344560 3732
rect 334676 3692 344560 3720
rect 334676 3680 334682 3692
rect 344554 3680 344560 3692
rect 344612 3680 344618 3732
rect 352834 3720 352840 3732
rect 344986 3692 352840 3720
rect 96338 3612 96344 3664
rect 96396 3652 96402 3664
rect 104526 3652 104532 3664
rect 96396 3624 104532 3652
rect 96396 3612 96402 3624
rect 104526 3612 104532 3624
rect 104584 3612 104590 3664
rect 107010 3612 107016 3664
rect 107068 3652 107074 3664
rect 115198 3652 115204 3664
rect 107068 3624 115204 3652
rect 107068 3612 107074 3624
rect 115198 3612 115204 3624
rect 115256 3612 115262 3664
rect 116670 3612 116676 3664
rect 116728 3652 116734 3664
rect 214650 3652 214656 3664
rect 116728 3624 214656 3652
rect 116728 3612 116734 3624
rect 214650 3612 214656 3624
rect 214708 3612 214714 3664
rect 224954 3612 224960 3664
rect 225012 3652 225018 3664
rect 277118 3652 277124 3664
rect 225012 3624 277124 3652
rect 225012 3612 225018 3624
rect 277118 3612 277124 3624
rect 277176 3612 277182 3664
rect 284294 3612 284300 3664
rect 284352 3652 284358 3664
rect 285030 3652 285036 3664
rect 284352 3624 285036 3652
rect 284352 3612 284358 3624
rect 285030 3612 285036 3624
rect 285088 3612 285094 3664
rect 285122 3612 285128 3664
rect 285180 3652 285186 3664
rect 304350 3652 304356 3664
rect 285180 3624 304356 3652
rect 285180 3612 285186 3624
rect 304350 3612 304356 3624
rect 304408 3612 304414 3664
rect 310422 3612 310428 3664
rect 310480 3652 310486 3664
rect 336274 3652 336280 3664
rect 310480 3624 336280 3652
rect 310480 3612 310486 3624
rect 336274 3612 336280 3624
rect 336332 3612 336338 3664
rect 340138 3612 340144 3664
rect 340196 3652 340202 3664
rect 344986 3652 345014 3692
rect 352834 3680 352840 3692
rect 352892 3680 352898 3732
rect 370958 3680 370964 3732
rect 371016 3720 371022 3732
rect 379974 3720 379980 3732
rect 371016 3692 379980 3720
rect 371016 3680 371022 3692
rect 379974 3680 379980 3692
rect 380032 3680 380038 3732
rect 389082 3680 389088 3732
rect 389140 3720 389146 3732
rect 394234 3720 394240 3732
rect 389140 3692 394240 3720
rect 389140 3680 389146 3692
rect 394234 3680 394240 3692
rect 394292 3680 394298 3732
rect 430574 3680 430580 3732
rect 430632 3720 430638 3732
rect 434438 3720 434444 3732
rect 430632 3692 434444 3720
rect 430632 3680 430638 3692
rect 434438 3680 434444 3692
rect 434496 3680 434502 3732
rect 448606 3680 448612 3732
rect 448664 3720 448670 3732
rect 514754 3720 514760 3732
rect 448664 3692 514760 3720
rect 448664 3680 448670 3692
rect 514754 3680 514760 3692
rect 514812 3680 514818 3732
rect 340196 3624 345014 3652
rect 340196 3612 340202 3624
rect 351914 3612 351920 3664
rect 351972 3652 351978 3664
rect 359918 3652 359924 3664
rect 351972 3624 359924 3652
rect 351972 3612 351978 3624
rect 359918 3612 359924 3624
rect 359976 3612 359982 3664
rect 377398 3612 377404 3664
rect 377456 3652 377462 3664
rect 388254 3652 388260 3664
rect 377456 3624 388260 3652
rect 377456 3612 377462 3624
rect 388254 3612 388260 3624
rect 388312 3612 388318 3664
rect 388438 3612 388444 3664
rect 388496 3652 388502 3664
rect 402514 3652 402520 3664
rect 388496 3624 402520 3652
rect 388496 3612 388502 3624
rect 402514 3612 402520 3624
rect 402572 3612 402578 3664
rect 403618 3612 403624 3664
rect 403676 3652 403682 3664
rect 420178 3652 420184 3664
rect 403676 3624 420184 3652
rect 403676 3612 403682 3624
rect 420178 3612 420184 3624
rect 420236 3612 420242 3664
rect 438762 3612 438768 3664
rect 438820 3652 438826 3664
rect 460382 3652 460388 3664
rect 438820 3624 460388 3652
rect 438820 3612 438826 3624
rect 460382 3612 460388 3624
rect 460440 3612 460446 3664
rect 462498 3612 462504 3664
rect 462556 3652 462562 3664
rect 533706 3652 533712 3664
rect 462556 3624 533712 3652
rect 462556 3612 462562 3624
rect 533706 3612 533712 3624
rect 533764 3612 533770 3664
rect 66956 3556 94452 3584
rect 66956 3544 66962 3556
rect 96890 3544 96896 3596
rect 96948 3584 96954 3596
rect 102226 3584 102232 3596
rect 96948 3556 102232 3584
rect 96948 3544 96954 3556
rect 102226 3544 102232 3556
rect 102284 3544 102290 3596
rect 102870 3544 102876 3596
rect 102928 3584 102934 3596
rect 103422 3584 103428 3596
rect 102928 3556 103428 3584
rect 102928 3544 102934 3556
rect 103422 3544 103428 3556
rect 103480 3544 103486 3596
rect 105078 3544 105084 3596
rect 105136 3584 105142 3596
rect 108482 3584 108488 3596
rect 105136 3556 108488 3584
rect 105136 3544 105142 3556
rect 108482 3544 108488 3556
rect 108540 3544 108546 3596
rect 108942 3544 108948 3596
rect 109000 3584 109006 3596
rect 109000 3556 109448 3584
rect 109000 3544 109006 3556
rect 81434 3516 81440 3528
rect 45526 3488 81440 3516
rect 81434 3476 81440 3488
rect 81492 3476 81498 3528
rect 88426 3476 88432 3528
rect 88484 3516 88490 3528
rect 108114 3516 108120 3528
rect 88484 3488 108120 3516
rect 88484 3476 88490 3488
rect 108114 3476 108120 3488
rect 108172 3476 108178 3528
rect 108298 3476 108304 3528
rect 108356 3516 108362 3528
rect 109310 3516 109316 3528
rect 108356 3488 109316 3516
rect 108356 3476 108362 3488
rect 109310 3476 109316 3488
rect 109368 3476 109374 3528
rect 109420 3516 109448 3556
rect 111058 3544 111064 3596
rect 111116 3584 111122 3596
rect 114002 3584 114008 3596
rect 111116 3556 114008 3584
rect 111116 3544 111122 3556
rect 114002 3544 114008 3556
rect 114060 3544 114066 3596
rect 117866 3544 117872 3596
rect 117924 3584 117930 3596
rect 433242 3584 433248 3596
rect 117924 3556 433248 3584
rect 117924 3544 117930 3556
rect 433242 3544 433248 3556
rect 433300 3544 433306 3596
rect 436002 3544 436008 3596
rect 436060 3584 436066 3596
rect 440326 3584 440332 3596
rect 436060 3556 440332 3584
rect 436060 3544 436066 3556
rect 440326 3544 440332 3556
rect 440384 3544 440390 3596
rect 440878 3544 440884 3596
rect 440936 3584 440942 3596
rect 452102 3584 452108 3596
rect 440936 3556 452108 3584
rect 440936 3544 440942 3556
rect 452102 3544 452108 3556
rect 452160 3544 452166 3596
rect 452746 3544 452752 3596
rect 452804 3584 452810 3596
rect 456886 3584 456892 3596
rect 452804 3556 456892 3584
rect 452804 3544 452810 3556
rect 456886 3544 456892 3556
rect 456944 3544 456950 3596
rect 457438 3544 457444 3596
rect 457496 3584 457502 3596
rect 537202 3584 537208 3596
rect 457496 3556 537208 3584
rect 457496 3544 457502 3556
rect 537202 3544 537208 3556
rect 537260 3544 537266 3596
rect 543734 3544 543740 3596
rect 543792 3584 543798 3596
rect 551462 3584 551468 3596
rect 543792 3556 551468 3584
rect 543792 3544 543798 3556
rect 551462 3544 551468 3556
rect 551520 3544 551526 3596
rect 116394 3516 116400 3528
rect 109420 3488 116400 3516
rect 116394 3476 116400 3488
rect 116452 3476 116458 3528
rect 118234 3476 118240 3528
rect 118292 3516 118298 3528
rect 468662 3516 468668 3528
rect 118292 3488 468668 3516
rect 118292 3476 118298 3488
rect 468662 3476 468668 3488
rect 468720 3476 468726 3528
rect 473814 3476 473820 3528
rect 473872 3516 473878 3528
rect 501782 3516 501788 3528
rect 473872 3488 501788 3516
rect 473872 3476 473878 3488
rect 501782 3476 501788 3488
rect 501840 3476 501846 3528
rect 503622 3476 503628 3528
rect 503680 3516 503686 3528
rect 505370 3516 505376 3528
rect 503680 3488 505376 3516
rect 503680 3476 503686 3488
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 509602 3476 509608 3528
rect 509660 3516 509666 3528
rect 523034 3516 523040 3528
rect 509660 3488 523040 3516
rect 509660 3476 509666 3488
rect 523034 3476 523040 3488
rect 523092 3476 523098 3528
rect 525794 3476 525800 3528
rect 525852 3516 525858 3528
rect 554958 3516 554964 3528
rect 525852 3488 554964 3516
rect 525852 3476 525858 3488
rect 554958 3476 554964 3488
rect 555016 3476 555022 3528
rect 562318 3476 562324 3528
rect 562376 3516 562382 3528
rect 564434 3516 564440 3528
rect 562376 3488 564440 3516
rect 562376 3476 562382 3488
rect 564434 3476 564440 3488
rect 564492 3476 564498 3528
rect 571242 3476 571248 3528
rect 571300 3516 571306 3528
rect 573910 3516 573916 3528
rect 571300 3488 573916 3516
rect 571300 3476 571306 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 17678 3448 17684 3460
rect 5316 3420 17684 3448
rect 5316 3408 5322 3420
rect 17678 3408 17684 3420
rect 17736 3408 17742 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 20680 3420 26234 3448
rect 20680 3408 20686 3420
rect 26206 3380 26234 3420
rect 40678 3408 40684 3460
rect 40736 3448 40742 3460
rect 43622 3448 43628 3460
rect 40736 3420 43628 3448
rect 40736 3408 40742 3420
rect 43622 3408 43628 3420
rect 43680 3408 43686 3460
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 47026 3448 47032 3460
rect 45520 3420 47032 3448
rect 45520 3408 45526 3420
rect 47026 3408 47032 3420
rect 47084 3408 47090 3460
rect 47486 3408 47492 3460
rect 47544 3448 47550 3460
rect 48958 3448 48964 3460
rect 47544 3420 48964 3448
rect 47544 3408 47550 3420
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 50338 3408 50344 3460
rect 50396 3448 50402 3460
rect 51350 3448 51356 3460
rect 50396 3420 51356 3448
rect 50396 3408 50402 3420
rect 51350 3408 51356 3420
rect 51408 3408 51414 3460
rect 54754 3408 54760 3460
rect 54812 3448 54818 3460
rect 56042 3448 56048 3460
rect 54812 3420 56048 3448
rect 54812 3408 54818 3420
rect 56042 3408 56048 3420
rect 56100 3408 56106 3460
rect 60090 3408 60096 3460
rect 60148 3448 60154 3460
rect 110506 3448 110512 3460
rect 60148 3420 110512 3448
rect 60148 3408 60154 3420
rect 110506 3408 110512 3420
rect 110564 3408 110570 3460
rect 113910 3408 113916 3460
rect 113968 3448 113974 3460
rect 475746 3448 475752 3460
rect 113968 3420 475752 3448
rect 113968 3408 113974 3420
rect 475746 3408 475752 3420
rect 475804 3408 475810 3460
rect 492030 3408 492036 3460
rect 492088 3448 492094 3460
rect 580994 3448 581000 3460
rect 492088 3420 581000 3448
rect 492088 3408 492094 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 42242 3380 42248 3392
rect 26206 3352 42248 3380
rect 42242 3340 42248 3352
rect 42300 3340 42306 3392
rect 50706 3340 50712 3392
rect 50764 3380 50770 3392
rect 54938 3380 54944 3392
rect 50764 3352 54944 3380
rect 50764 3340 50770 3352
rect 54938 3340 54944 3352
rect 54996 3340 55002 3392
rect 59630 3380 59636 3392
rect 55186 3352 59636 3380
rect 35986 3272 35992 3324
rect 36044 3312 36050 3324
rect 39298 3312 39304 3324
rect 36044 3284 39304 3312
rect 36044 3272 36050 3284
rect 39298 3272 39304 3284
rect 39356 3272 39362 3324
rect 49142 3272 49148 3324
rect 49200 3312 49206 3324
rect 55186 3312 55214 3352
rect 59630 3340 59636 3352
rect 59688 3340 59694 3392
rect 79502 3340 79508 3392
rect 79560 3380 79566 3392
rect 98638 3380 98644 3392
rect 79560 3352 98644 3380
rect 79560 3340 79566 3352
rect 98638 3340 98644 3352
rect 98696 3340 98702 3392
rect 99834 3380 99840 3392
rect 99346 3352 99840 3380
rect 49200 3284 55214 3312
rect 49200 3272 49206 3284
rect 84930 3272 84936 3324
rect 84988 3312 84994 3324
rect 91554 3312 91560 3324
rect 84988 3284 91560 3312
rect 84988 3272 84994 3284
rect 91554 3272 91560 3284
rect 91612 3272 91618 3324
rect 92934 3272 92940 3324
rect 92992 3312 92998 3324
rect 96246 3312 96252 3324
rect 92992 3284 96252 3312
rect 92992 3272 92998 3284
rect 96246 3272 96252 3284
rect 96304 3272 96310 3324
rect 97258 3272 97264 3324
rect 97316 3312 97322 3324
rect 99346 3312 99374 3352
rect 99834 3340 99840 3352
rect 99892 3340 99898 3392
rect 104802 3380 104808 3392
rect 99944 3352 104808 3380
rect 97316 3284 99374 3312
rect 97316 3272 97322 3284
rect 59998 3204 60004 3256
rect 60056 3244 60062 3256
rect 63218 3244 63224 3256
rect 60056 3216 63224 3244
rect 60056 3204 60062 3216
rect 63218 3204 63224 3216
rect 63276 3204 63282 3256
rect 82170 3204 82176 3256
rect 82228 3244 82234 3256
rect 95142 3244 95148 3256
rect 82228 3216 95148 3244
rect 82228 3204 82234 3216
rect 95142 3204 95148 3216
rect 95200 3204 95206 3256
rect 97994 3204 98000 3256
rect 98052 3244 98058 3256
rect 99944 3244 99972 3352
rect 104802 3340 104808 3352
rect 104860 3340 104866 3392
rect 108206 3340 108212 3392
rect 108264 3380 108270 3392
rect 121086 3380 121092 3392
rect 108264 3352 121092 3380
rect 108264 3340 108270 3352
rect 121086 3340 121092 3352
rect 121144 3340 121150 3392
rect 121270 3340 121276 3392
rect 121328 3380 121334 3392
rect 128170 3380 128176 3392
rect 121328 3352 128176 3380
rect 121328 3340 121334 3352
rect 128170 3340 128176 3352
rect 128228 3340 128234 3392
rect 131206 3340 131212 3392
rect 131264 3380 131270 3392
rect 135254 3380 135260 3392
rect 131264 3352 135260 3380
rect 131264 3340 131270 3352
rect 135254 3340 135260 3352
rect 135312 3340 135318 3392
rect 149514 3340 149520 3392
rect 149572 3380 149578 3392
rect 151354 3380 151360 3392
rect 149572 3352 151360 3380
rect 149572 3340 149578 3352
rect 151354 3340 151360 3352
rect 151412 3340 151418 3392
rect 155402 3380 155408 3392
rect 151786 3352 155408 3380
rect 111610 3312 111616 3324
rect 98052 3216 99972 3244
rect 100036 3284 111616 3312
rect 98052 3204 98058 3216
rect 39574 3136 39580 3188
rect 39632 3176 39638 3188
rect 42058 3176 42064 3188
rect 39632 3148 42064 3176
rect 39632 3136 39638 3148
rect 42058 3136 42064 3148
rect 42116 3136 42122 3188
rect 92382 3136 92388 3188
rect 92440 3176 92446 3188
rect 100036 3176 100064 3284
rect 111610 3272 111616 3284
rect 111668 3272 111674 3324
rect 111794 3272 111800 3324
rect 111852 3312 111858 3324
rect 117866 3312 117872 3324
rect 111852 3284 117872 3312
rect 111852 3272 111858 3284
rect 117866 3272 117872 3284
rect 117924 3272 117930 3324
rect 146662 3272 146668 3324
rect 146720 3312 146726 3324
rect 151786 3312 151814 3352
rect 155402 3340 155408 3352
rect 155460 3340 155466 3392
rect 160094 3340 160100 3392
rect 160152 3380 160158 3392
rect 161290 3380 161296 3392
rect 160152 3352 161296 3380
rect 160152 3340 160158 3352
rect 161290 3340 161296 3352
rect 161348 3340 161354 3392
rect 174538 3340 174544 3392
rect 174596 3380 174602 3392
rect 176654 3380 176660 3392
rect 174596 3352 176660 3380
rect 174596 3340 174602 3352
rect 176654 3340 176660 3352
rect 176712 3340 176718 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186130 3380 186136 3392
rect 184992 3352 186136 3380
rect 184992 3340 184998 3352
rect 186130 3340 186136 3352
rect 186188 3340 186194 3392
rect 299474 3340 299480 3392
rect 299532 3380 299538 3392
rect 300762 3380 300768 3392
rect 299532 3352 300768 3380
rect 299532 3340 299538 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 307846 3340 307852 3392
rect 307904 3380 307910 3392
rect 309042 3380 309048 3392
rect 307904 3352 309048 3380
rect 307904 3340 307910 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 354674 3340 354680 3392
rect 354732 3380 354738 3392
rect 358722 3380 358728 3392
rect 354732 3352 358728 3380
rect 354732 3340 354738 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 358814 3340 358820 3392
rect 358872 3380 358878 3392
rect 362310 3380 362316 3392
rect 358872 3352 362316 3380
rect 358872 3340 358878 3352
rect 362310 3340 362316 3352
rect 362368 3340 362374 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 146720 3284 151814 3312
rect 146720 3272 146726 3284
rect 160554 3272 160560 3324
rect 160612 3312 160618 3324
rect 163682 3312 163688 3324
rect 160612 3284 163688 3312
rect 160612 3272 160618 3284
rect 163682 3272 163688 3284
rect 163740 3272 163746 3324
rect 223482 3272 223488 3324
rect 223540 3312 223546 3324
rect 231026 3312 231032 3324
rect 223540 3284 231032 3312
rect 223540 3272 223546 3284
rect 231026 3272 231032 3284
rect 231084 3272 231090 3324
rect 252462 3272 252468 3324
rect 252520 3312 252526 3324
rect 259454 3312 259460 3324
rect 252520 3284 259460 3312
rect 252520 3272 252526 3284
rect 259454 3272 259460 3284
rect 259512 3272 259518 3324
rect 321462 3272 321468 3324
rect 321520 3312 321526 3324
rect 323302 3312 323308 3324
rect 321520 3284 323308 3312
rect 321520 3272 321526 3284
rect 323302 3272 323308 3284
rect 323360 3272 323366 3324
rect 372614 3272 372620 3324
rect 372672 3312 372678 3324
rect 376478 3312 376484 3324
rect 372672 3284 376484 3312
rect 372672 3272 372678 3284
rect 376478 3272 376484 3284
rect 376536 3272 376542 3324
rect 484394 3272 484400 3324
rect 484452 3312 484458 3324
rect 487614 3312 487620 3324
rect 484452 3284 487620 3312
rect 484452 3272 484458 3284
rect 487614 3272 487620 3284
rect 487672 3272 487678 3324
rect 565814 3272 565820 3324
rect 565872 3312 565878 3324
rect 569126 3312 569132 3324
rect 565872 3284 569132 3312
rect 565872 3272 565878 3284
rect 569126 3272 569132 3284
rect 569184 3272 569190 3324
rect 101306 3204 101312 3256
rect 101364 3244 101370 3256
rect 118786 3244 118792 3256
rect 101364 3216 118792 3244
rect 101364 3204 101370 3216
rect 118786 3204 118792 3216
rect 118844 3204 118850 3256
rect 471882 3204 471888 3256
rect 471940 3244 471946 3256
rect 473446 3244 473452 3256
rect 471940 3216 473452 3244
rect 471940 3204 471946 3216
rect 473446 3204 473452 3216
rect 473504 3204 473510 3256
rect 92440 3148 100064 3176
rect 92440 3136 92446 3148
rect 102594 3136 102600 3188
rect 102652 3176 102658 3188
rect 117590 3176 117596 3188
rect 102652 3148 117596 3176
rect 102652 3136 102658 3148
rect 117590 3136 117596 3148
rect 117648 3136 117654 3188
rect 124582 3136 124588 3188
rect 124640 3176 124646 3188
rect 156966 3176 156972 3188
rect 124640 3148 156972 3176
rect 124640 3136 124646 3148
rect 156966 3136 156972 3148
rect 157024 3136 157030 3188
rect 162854 3136 162860 3188
rect 162912 3176 162918 3188
rect 169570 3176 169576 3188
rect 162912 3148 169576 3176
rect 162912 3136 162918 3148
rect 169570 3136 169576 3148
rect 169628 3136 169634 3188
rect 221642 3136 221648 3188
rect 221700 3176 221706 3188
rect 223942 3176 223948 3188
rect 221700 3148 223948 3176
rect 221700 3136 221706 3148
rect 223942 3136 223948 3148
rect 224000 3136 224006 3188
rect 360102 3136 360108 3188
rect 360160 3176 360166 3188
rect 363506 3176 363512 3188
rect 360160 3148 363512 3176
rect 360160 3136 360166 3148
rect 363506 3136 363512 3148
rect 363564 3136 363570 3188
rect 413278 3136 413284 3188
rect 413336 3176 413342 3188
rect 416682 3176 416688 3188
rect 413336 3148 416688 3176
rect 413336 3136 413342 3148
rect 416682 3136 416688 3148
rect 416740 3136 416746 3188
rect 434622 3136 434628 3188
rect 434680 3176 434686 3188
rect 437934 3176 437940 3188
rect 434680 3148 437940 3176
rect 434680 3136 434686 3148
rect 437934 3136 437940 3148
rect 437992 3136 437998 3188
rect 481542 3136 481548 3188
rect 481600 3176 481606 3188
rect 484026 3176 484032 3188
rect 481600 3148 484032 3176
rect 481600 3136 481606 3148
rect 484026 3136 484032 3148
rect 484084 3136 484090 3188
rect 512638 3136 512644 3188
rect 512696 3176 512702 3188
rect 515950 3176 515956 3188
rect 512696 3148 515956 3176
rect 512696 3136 512702 3148
rect 515950 3136 515956 3148
rect 516008 3136 516014 3188
rect 91738 3068 91744 3120
rect 91796 3108 91802 3120
rect 105722 3108 105728 3120
rect 91796 3080 105728 3108
rect 91796 3068 91802 3080
rect 105722 3068 105728 3080
rect 105780 3068 105786 3120
rect 191742 3068 191748 3120
rect 191800 3108 191806 3120
rect 195606 3108 195612 3120
rect 191800 3080 195612 3108
rect 191800 3068 191806 3080
rect 195606 3068 195612 3080
rect 195664 3068 195670 3120
rect 220722 3068 220728 3120
rect 220780 3108 220786 3120
rect 246390 3108 246396 3120
rect 220780 3080 246396 3108
rect 220780 3068 220786 3080
rect 246390 3068 246396 3080
rect 246448 3068 246454 3120
rect 291838 3068 291844 3120
rect 291896 3108 291902 3120
rect 294874 3108 294880 3120
rect 291896 3080 294880 3108
rect 291896 3068 291902 3080
rect 294874 3068 294880 3080
rect 294932 3068 294938 3120
rect 294966 3068 294972 3120
rect 295024 3108 295030 3120
rect 298462 3108 298468 3120
rect 295024 3080 298468 3108
rect 295024 3068 295030 3080
rect 298462 3068 298468 3080
rect 298520 3068 298526 3120
rect 445110 3068 445116 3120
rect 445168 3108 445174 3120
rect 448606 3108 448612 3120
rect 445168 3080 448612 3108
rect 445168 3068 445174 3080
rect 448606 3068 448612 3080
rect 448664 3068 448670 3120
rect 103974 3000 103980 3052
rect 104032 3040 104038 3052
rect 108574 3040 108580 3052
rect 104032 3012 108580 3040
rect 104032 3000 104038 3012
rect 108574 3000 108580 3012
rect 108632 3000 108638 3052
rect 150434 3000 150440 3052
rect 150492 3040 150498 3052
rect 153838 3040 153844 3052
rect 150492 3012 153844 3040
rect 150492 3000 150498 3012
rect 153838 3000 153844 3012
rect 153896 3000 153902 3052
rect 157334 3000 157340 3052
rect 157392 3040 157398 3052
rect 232222 3040 232228 3052
rect 157392 3012 232228 3040
rect 157392 3000 157398 3012
rect 232222 3000 232228 3012
rect 232280 3000 232286 3052
rect 278038 3000 278044 3052
rect 278096 3040 278102 3052
rect 280706 3040 280712 3052
rect 278096 3012 280712 3040
rect 278096 3000 278102 3012
rect 280706 3000 280712 3012
rect 280764 3000 280770 3052
rect 395430 3000 395436 3052
rect 395488 3040 395494 3052
rect 397730 3040 397736 3052
rect 395488 3012 397736 3040
rect 395488 3000 395494 3012
rect 397730 3000 397736 3012
rect 397788 3000 397794 3052
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 3418 2972 3424 2984
rect 1728 2944 3424 2972
rect 1728 2932 1734 2944
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 37182 2932 37188 2984
rect 37240 2972 37246 2984
rect 43530 2972 43536 2984
rect 37240 2944 43536 2972
rect 37240 2932 37246 2944
rect 43530 2932 43536 2944
rect 43588 2932 43594 2984
rect 133782 2932 133788 2984
rect 133840 2972 133846 2984
rect 138842 2972 138848 2984
rect 133840 2944 138848 2972
rect 133840 2932 133846 2944
rect 138842 2932 138848 2944
rect 138900 2932 138906 2984
rect 139394 2932 139400 2984
rect 139452 2972 139458 2984
rect 142430 2972 142436 2984
rect 139452 2944 142436 2972
rect 139452 2932 139458 2944
rect 142430 2932 142436 2944
rect 142488 2932 142494 2984
rect 194962 2932 194968 2984
rect 195020 2972 195026 2984
rect 214466 2972 214472 2984
rect 195020 2944 214472 2972
rect 195020 2932 195026 2944
rect 214466 2932 214472 2944
rect 214524 2932 214530 2984
rect 214558 2932 214564 2984
rect 214616 2972 214622 2984
rect 235810 2972 235816 2984
rect 214616 2944 235816 2972
rect 214616 2932 214622 2944
rect 235810 2932 235816 2944
rect 235868 2932 235874 2984
rect 322198 2932 322204 2984
rect 322256 2972 322262 2984
rect 326798 2972 326804 2984
rect 322256 2944 326804 2972
rect 322256 2932 322262 2944
rect 326798 2932 326804 2944
rect 326856 2932 326862 2984
rect 118602 2864 118608 2916
rect 118660 2904 118666 2916
rect 122282 2904 122288 2916
rect 118660 2876 122288 2904
rect 118660 2864 118666 2876
rect 122282 2864 122288 2876
rect 122340 2864 122346 2916
rect 129734 2864 129740 2916
rect 129792 2904 129798 2916
rect 141234 2904 141240 2916
rect 129792 2876 141240 2904
rect 129792 2864 129798 2876
rect 141234 2864 141240 2876
rect 141292 2864 141298 2916
rect 154482 2864 154488 2916
rect 154540 2904 154546 2916
rect 157794 2904 157800 2916
rect 154540 2876 157800 2904
rect 154540 2864 154546 2876
rect 157794 2864 157800 2876
rect 157852 2864 157858 2916
rect 201034 2864 201040 2916
rect 201092 2904 201098 2916
rect 221550 2904 221556 2916
rect 201092 2876 221556 2904
rect 201092 2864 201098 2876
rect 221550 2864 221556 2876
rect 221608 2864 221614 2916
rect 258718 2864 258724 2916
rect 258776 2904 258782 2916
rect 262950 2904 262956 2916
rect 258776 2876 262956 2904
rect 258776 2864 258782 2876
rect 262950 2864 262956 2876
rect 263008 2864 263014 2916
rect 363046 2864 363052 2916
rect 363104 2904 363110 2916
rect 365806 2904 365812 2916
rect 363104 2876 365812 2904
rect 363104 2864 363110 2876
rect 365806 2864 365812 2876
rect 365864 2864 365870 2916
rect 368382 2864 368388 2916
rect 368440 2904 368446 2916
rect 370590 2904 370596 2916
rect 368440 2876 370596 2904
rect 368440 2864 368446 2876
rect 370590 2864 370596 2876
rect 370648 2864 370654 2916
rect 115842 2796 115848 2848
rect 115900 2836 115906 2848
rect 144730 2836 144736 2848
rect 115900 2808 117360 2836
rect 115900 2796 115906 2808
rect 33134 2728 33140 2780
rect 33192 2768 33198 2780
rect 112162 2768 112168 2780
rect 33192 2740 112168 2768
rect 33192 2728 33198 2740
rect 112162 2728 112168 2740
rect 112220 2728 112226 2780
rect 112438 2728 112444 2780
rect 112496 2768 112502 2780
rect 114462 2768 114468 2780
rect 112496 2740 114468 2768
rect 112496 2728 112502 2740
rect 114462 2728 114468 2740
rect 114520 2728 114526 2780
rect 117332 2768 117360 2808
rect 120092 2808 129780 2836
rect 120092 2768 120120 2808
rect 117332 2740 120120 2768
rect 129752 2768 129780 2808
rect 136560 2808 144736 2836
rect 136560 2768 136588 2808
rect 144730 2796 144736 2808
rect 144788 2796 144794 2848
rect 153010 2796 153016 2848
rect 153068 2836 153074 2848
rect 158898 2836 158904 2848
rect 153068 2808 158904 2836
rect 153068 2796 153074 2808
rect 158898 2796 158904 2808
rect 158956 2796 158962 2848
rect 202782 2796 202788 2848
rect 202840 2836 202846 2848
rect 208578 2836 208584 2848
rect 202840 2808 208584 2836
rect 202840 2796 202846 2808
rect 208578 2796 208584 2808
rect 208636 2796 208642 2848
rect 218146 2796 218152 2848
rect 218204 2836 218210 2848
rect 225138 2836 225144 2848
rect 218204 2808 225144 2836
rect 218204 2796 218210 2808
rect 225138 2796 225144 2808
rect 225196 2796 225202 2848
rect 247034 2796 247040 2848
rect 247092 2836 247098 2848
rect 249978 2836 249984 2848
rect 247092 2808 249984 2836
rect 247092 2796 247098 2808
rect 249978 2796 249984 2808
rect 250036 2796 250042 2848
rect 274634 2796 274640 2848
rect 274692 2836 274698 2848
rect 279510 2836 279516 2848
rect 274692 2808 279516 2836
rect 274692 2796 274698 2808
rect 279510 2796 279516 2808
rect 279568 2796 279574 2848
rect 409782 2796 409788 2848
rect 409840 2836 409846 2848
rect 411898 2836 411904 2848
rect 409840 2808 411904 2836
rect 409840 2796 409846 2808
rect 411898 2796 411904 2808
rect 411956 2796 411962 2848
rect 427722 2796 427728 2848
rect 427780 2836 427786 2848
rect 429654 2836 429660 2848
rect 427780 2808 429660 2836
rect 427780 2796 427786 2808
rect 429654 2796 429660 2808
rect 429712 2796 429718 2848
rect 445662 2796 445668 2848
rect 445720 2836 445726 2848
rect 447410 2836 447416 2848
rect 445720 2808 447416 2836
rect 445720 2796 445726 2808
rect 447410 2796 447416 2808
rect 447468 2796 447474 2848
rect 521562 2796 521568 2848
rect 521620 2836 521626 2848
rect 524230 2836 524236 2848
rect 521620 2808 524236 2836
rect 521620 2796 521626 2808
rect 524230 2796 524236 2808
rect 524288 2796 524294 2848
rect 552566 2796 552572 2848
rect 552624 2836 552630 2848
rect 559742 2836 559748 2848
rect 552624 2808 559748 2836
rect 552624 2796 552630 2808
rect 559742 2796 559748 2808
rect 559800 2796 559806 2848
rect 572714 2836 572720 2848
rect 571260 2808 572720 2836
rect 129752 2740 136588 2768
rect 149606 2728 149612 2780
rect 149664 2768 149670 2780
rect 571260 2768 571288 2808
rect 572714 2796 572720 2808
rect 572772 2796 572778 2848
rect 149664 2740 571288 2768
rect 149664 2728 149670 2740
rect 76558 2660 76564 2712
rect 76616 2700 76622 2712
rect 214558 2700 214564 2712
rect 76616 2672 214564 2700
rect 76616 2660 76622 2672
rect 214558 2660 214564 2672
rect 214616 2660 214622 2712
rect 214650 2660 214656 2712
rect 214708 2700 214714 2712
rect 445662 2700 445668 2712
rect 214708 2672 445668 2700
rect 214708 2660 214714 2672
rect 445662 2660 445668 2672
rect 445720 2660 445726 2712
rect 116578 2592 116584 2644
rect 116636 2632 116642 2644
rect 117866 2632 117872 2644
rect 116636 2604 117872 2632
rect 116636 2592 116642 2604
rect 117866 2592 117872 2604
rect 117924 2592 117930 2644
rect 124214 2592 124220 2644
rect 124272 2632 124278 2644
rect 130562 2632 130568 2644
rect 124272 2604 130568 2632
rect 124272 2592 124278 2604
rect 130562 2592 130568 2604
rect 130620 2592 130626 2644
rect 143902 2592 143908 2644
rect 143960 2632 143966 2644
rect 153746 2632 153752 2644
rect 143960 2604 153752 2632
rect 143960 2592 143966 2604
rect 153746 2592 153752 2604
rect 153804 2592 153810 2644
rect 195974 2592 195980 2644
rect 196032 2632 196038 2644
rect 409782 2632 409788 2644
rect 196032 2604 409788 2632
rect 196032 2592 196038 2604
rect 409782 2592 409788 2604
rect 409840 2592 409846 2644
rect 78214 2524 78220 2576
rect 78272 2564 78278 2576
rect 220722 2564 220728 2576
rect 78272 2536 220728 2564
rect 78272 2524 78278 2536
rect 220722 2524 220728 2536
rect 220780 2524 220786 2576
rect 58894 2456 58900 2508
rect 58952 2496 58958 2508
rect 118602 2496 118608 2508
rect 58952 2468 118608 2496
rect 58952 2456 58958 2468
rect 118602 2456 118608 2468
rect 118660 2456 118666 2508
rect 157334 2496 157340 2508
rect 128326 2468 157340 2496
rect 76006 2388 76012 2440
rect 76064 2428 76070 2440
rect 128326 2428 128354 2468
rect 157334 2456 157340 2468
rect 157392 2456 157398 2508
rect 173526 2456 173532 2508
rect 173584 2496 173590 2508
rect 202782 2496 202788 2508
rect 173584 2468 202788 2496
rect 173584 2456 173590 2468
rect 202782 2456 202788 2468
rect 202840 2456 202846 2508
rect 76064 2400 128354 2428
rect 76064 2388 76070 2400
rect 158806 2388 158812 2440
rect 158864 2428 158870 2440
rect 218146 2428 218152 2440
rect 158864 2400 218152 2428
rect 158864 2388 158870 2400
rect 218146 2388 218152 2400
rect 218204 2388 218210 2440
rect 237374 2388 237380 2440
rect 237432 2428 237438 2440
rect 247034 2428 247040 2440
rect 237432 2400 247040 2428
rect 237432 2388 237438 2400
rect 247034 2388 247040 2400
rect 247092 2388 247098 2440
rect 67910 2320 67916 2372
rect 67968 2360 67974 2372
rect 112070 2360 112076 2372
rect 67968 2332 112076 2360
rect 67968 2320 67974 2332
rect 112070 2320 112076 2332
rect 112128 2320 112134 2372
rect 120718 2320 120724 2372
rect 120776 2360 120782 2372
rect 274818 2360 274824 2372
rect 120776 2332 274824 2360
rect 120776 2320 120782 2332
rect 274818 2320 274824 2332
rect 274876 2320 274882 2372
rect 87598 2252 87604 2304
rect 87656 2292 87662 2304
rect 264146 2292 264152 2304
rect 87656 2264 264152 2292
rect 87656 2252 87662 2264
rect 264146 2252 264152 2264
rect 264204 2252 264210 2304
rect 81434 2184 81440 2236
rect 81492 2224 81498 2236
rect 87138 2224 87144 2236
rect 81492 2196 87144 2224
rect 81492 2184 81498 2196
rect 87138 2184 87144 2196
rect 87196 2184 87202 2236
rect 91646 2184 91652 2236
rect 91704 2224 91710 2236
rect 278314 2224 278320 2236
rect 91704 2196 278320 2224
rect 91704 2184 91710 2196
rect 278314 2184 278320 2196
rect 278372 2184 278378 2236
rect 60734 2116 60740 2168
rect 60792 2156 60798 2168
rect 132954 2156 132960 2168
rect 60792 2128 132960 2156
rect 60792 2116 60798 2128
rect 132954 2116 132960 2128
rect 133012 2116 133018 2168
rect 135070 2116 135076 2168
rect 135128 2156 135134 2168
rect 144822 2156 144828 2168
rect 135128 2128 144828 2156
rect 135128 2116 135134 2128
rect 144822 2116 144828 2128
rect 144880 2116 144886 2168
rect 144914 2116 144920 2168
rect 144972 2156 144978 2168
rect 194962 2156 194968 2168
rect 144972 2128 194968 2156
rect 144972 2116 144978 2128
rect 194962 2116 194968 2128
rect 195020 2116 195026 2168
rect 200666 2116 200672 2168
rect 200724 2156 200730 2168
rect 404814 2156 404820 2168
rect 200724 2128 404820 2156
rect 200724 2116 200730 2128
rect 404814 2116 404820 2128
rect 404872 2116 404878 2168
rect 63494 2048 63500 2100
rect 63552 2088 63558 2100
rect 63552 2060 138014 2088
rect 63552 2048 63558 2060
rect 74350 1980 74356 2032
rect 74408 2020 74414 2032
rect 106182 2020 106188 2032
rect 74408 1992 106188 2020
rect 74408 1980 74414 1992
rect 106182 1980 106188 1992
rect 106240 1980 106246 2032
rect 112530 1980 112536 2032
rect 112588 2020 112594 2032
rect 129734 2020 129740 2032
rect 112588 1992 129740 2020
rect 112588 1980 112594 1992
rect 129734 1980 129740 1992
rect 129792 1980 129798 2032
rect 75454 1912 75460 1964
rect 75512 1952 75518 1964
rect 100754 1952 100760 1964
rect 75512 1924 100760 1952
rect 75512 1912 75518 1924
rect 100754 1912 100760 1924
rect 100812 1912 100818 1964
rect 104802 1912 104808 1964
rect 104860 1952 104866 1964
rect 121454 1952 121460 1964
rect 104860 1924 121460 1952
rect 104860 1912 104866 1924
rect 121454 1912 121460 1924
rect 121512 1912 121518 1964
rect 137986 1952 138014 2060
rect 153102 2048 153108 2100
rect 153160 2088 153166 2100
rect 201034 2088 201040 2100
rect 153160 2060 201040 2088
rect 153160 2048 153166 2060
rect 201034 2048 201040 2060
rect 201092 2048 201098 2100
rect 201678 2048 201684 2100
rect 201736 2088 201742 2100
rect 418982 2088 418988 2100
rect 201736 2060 418988 2088
rect 201736 2048 201742 2060
rect 418982 2048 418988 2060
rect 419040 2048 419046 2100
rect 140774 1980 140780 2032
rect 140832 2020 140838 2032
rect 154482 2020 154488 2032
rect 140832 1992 154488 2020
rect 140832 1980 140838 1992
rect 154482 1980 154488 1992
rect 154540 1980 154546 2032
rect 151814 1952 151820 1964
rect 137986 1924 151820 1952
rect 151814 1912 151820 1924
rect 151872 1912 151878 1964
rect 97534 1844 97540 1896
rect 97592 1884 97598 1896
rect 115842 1884 115848 1896
rect 97592 1856 115848 1884
rect 97592 1844 97598 1856
rect 115842 1844 115848 1856
rect 115900 1844 115906 1896
rect 80698 1776 80704 1828
rect 80756 1816 80762 1828
rect 150434 1816 150440 1828
rect 80756 1788 150440 1816
rect 80756 1776 80762 1788
rect 150434 1776 150440 1788
rect 150492 1776 150498 1828
rect 121178 1640 121184 1692
rect 121236 1680 121242 1692
rect 124122 1680 124128 1692
rect 121236 1652 124128 1680
rect 121236 1640 121242 1652
rect 124122 1640 124128 1652
rect 124180 1640 124186 1692
rect 137278 1640 137284 1692
rect 137336 1680 137342 1692
rect 178034 1680 178040 1692
rect 137336 1652 178040 1680
rect 137336 1640 137342 1652
rect 178034 1640 178040 1652
rect 178092 1640 178098 1692
rect 121362 1572 121368 1624
rect 121420 1612 121426 1624
rect 128354 1612 128360 1624
rect 121420 1584 128360 1612
rect 121420 1572 121426 1584
rect 128354 1572 128360 1584
rect 128412 1572 128418 1624
rect 142798 1612 142804 1624
rect 132466 1584 142804 1612
rect 122834 1504 122840 1556
rect 122892 1544 122898 1556
rect 124858 1544 124864 1556
rect 122892 1516 124864 1544
rect 122892 1504 122898 1516
rect 124858 1504 124864 1516
rect 124916 1504 124922 1556
rect 122742 1436 122748 1488
rect 122800 1476 122806 1488
rect 125870 1476 125876 1488
rect 122800 1448 125876 1476
rect 122800 1436 122806 1448
rect 125870 1436 125876 1448
rect 125928 1436 125934 1488
rect 132466 1476 132494 1584
rect 142798 1572 142804 1584
rect 142856 1572 142862 1624
rect 136542 1504 136548 1556
rect 136600 1544 136606 1556
rect 146294 1544 146300 1556
rect 136600 1516 146300 1544
rect 136600 1504 136606 1516
rect 146294 1504 146300 1516
rect 146352 1504 146358 1556
rect 128326 1448 132494 1476
rect 122926 1408 122932 1420
rect 103486 1380 122932 1408
rect 85942 1232 85948 1284
rect 86000 1272 86006 1284
rect 103486 1272 103514 1380
rect 122926 1368 122932 1380
rect 122984 1368 122990 1420
rect 123018 1368 123024 1420
rect 123076 1408 123082 1420
rect 128326 1408 128354 1448
rect 133782 1436 133788 1488
rect 133840 1476 133846 1488
rect 140038 1476 140044 1488
rect 133840 1448 140044 1476
rect 133840 1436 133846 1448
rect 140038 1436 140044 1448
rect 140096 1436 140102 1488
rect 149054 1476 149060 1488
rect 142816 1448 149060 1476
rect 123076 1380 128354 1408
rect 129752 1380 135208 1408
rect 123076 1368 123082 1380
rect 115842 1300 115848 1352
rect 115900 1340 115906 1352
rect 121178 1340 121184 1352
rect 115900 1312 121184 1340
rect 115900 1300 115906 1312
rect 121178 1300 121184 1312
rect 121236 1300 121242 1352
rect 126974 1300 126980 1352
rect 127032 1340 127038 1352
rect 129752 1340 129780 1380
rect 127032 1312 129780 1340
rect 135180 1340 135208 1380
rect 136266 1368 136272 1420
rect 136324 1408 136330 1420
rect 142816 1408 142844 1448
rect 149054 1436 149060 1448
rect 149112 1436 149118 1488
rect 218238 1436 218244 1488
rect 218296 1476 218302 1488
rect 228726 1476 228732 1488
rect 218296 1448 228732 1476
rect 218296 1436 218302 1448
rect 228726 1436 228732 1448
rect 228784 1436 228790 1488
rect 136324 1380 142844 1408
rect 136324 1368 136330 1380
rect 142890 1368 142896 1420
rect 142948 1408 142954 1420
rect 158714 1408 158720 1420
rect 142948 1380 144960 1408
rect 142948 1368 142954 1380
rect 137278 1340 137284 1352
rect 135180 1312 137284 1340
rect 127032 1300 127038 1312
rect 137278 1300 137284 1312
rect 137336 1300 137342 1352
rect 144932 1340 144960 1380
rect 147692 1380 158720 1408
rect 147692 1340 147720 1380
rect 158714 1368 158720 1380
rect 158772 1368 158778 1420
rect 239306 1408 239312 1420
rect 178052 1380 239312 1408
rect 144932 1312 147720 1340
rect 148318 1300 148324 1352
rect 148376 1340 148382 1352
rect 150802 1340 150808 1352
rect 148376 1312 150808 1340
rect 148376 1300 148382 1312
rect 150802 1300 150808 1312
rect 150860 1300 150866 1352
rect 86000 1244 103514 1272
rect 86000 1232 86006 1244
rect 114462 1232 114468 1284
rect 114520 1272 114526 1284
rect 121362 1272 121368 1284
rect 114520 1244 121368 1272
rect 114520 1232 114526 1244
rect 121362 1232 121368 1244
rect 121420 1232 121426 1284
rect 121454 1232 121460 1284
rect 121512 1272 121518 1284
rect 129642 1272 129648 1284
rect 121512 1244 129648 1272
rect 121512 1232 121518 1244
rect 129642 1232 129648 1244
rect 129700 1232 129706 1284
rect 146294 1232 146300 1284
rect 146352 1272 146358 1284
rect 149238 1272 149244 1284
rect 146352 1244 149244 1272
rect 146352 1232 146358 1244
rect 149238 1232 149244 1244
rect 149296 1232 149302 1284
rect 64874 1164 64880 1216
rect 64932 1204 64938 1216
rect 114094 1204 114100 1216
rect 64932 1176 114100 1204
rect 64932 1164 64938 1176
rect 114094 1164 114100 1176
rect 114152 1164 114158 1216
rect 139486 1164 139492 1216
rect 139544 1204 139550 1216
rect 153010 1204 153016 1216
rect 139544 1176 153016 1204
rect 139544 1164 139550 1176
rect 153010 1164 153016 1176
rect 153068 1164 153074 1216
rect 77110 1096 77116 1148
rect 77168 1136 77174 1148
rect 178052 1136 178080 1380
rect 239306 1368 239312 1380
rect 239364 1368 239370 1420
rect 276014 1368 276020 1420
rect 276072 1408 276078 1420
rect 281902 1408 281908 1420
rect 276072 1380 281908 1408
rect 276072 1368 276078 1380
rect 281902 1368 281908 1380
rect 281960 1368 281966 1420
rect 313274 1368 313280 1420
rect 313332 1408 313338 1420
rect 320910 1408 320916 1420
rect 313332 1380 320916 1408
rect 313332 1368 313338 1380
rect 320910 1368 320916 1380
rect 320968 1368 320974 1420
rect 77168 1108 178080 1136
rect 77168 1096 77174 1108
rect 72326 1028 72332 1080
rect 72384 1068 72390 1080
rect 173526 1068 173532 1080
rect 72384 1040 173532 1068
rect 72384 1028 72390 1040
rect 173526 1028 173532 1040
rect 173584 1028 173590 1080
rect 69658 960 69664 1012
rect 69716 1000 69722 1012
rect 133782 1000 133788 1012
rect 69716 972 133788 1000
rect 69716 960 69722 972
rect 133782 960 133788 972
rect 133840 960 133846 1012
rect 142798 960 142804 1012
rect 142856 1000 142862 1012
rect 158806 1000 158812 1012
rect 142856 972 158812 1000
rect 142856 960 142862 972
rect 158806 960 158812 972
rect 158864 960 158870 1012
rect 60918 892 60924 944
rect 60976 932 60982 944
rect 122742 932 122748 944
rect 60976 904 122748 932
rect 60976 892 60982 904
rect 122742 892 122748 904
rect 122800 892 122806 944
rect 122926 892 122932 944
rect 122984 932 122990 944
rect 142890 932 142896 944
rect 122984 904 142896 932
rect 122984 892 122990 904
rect 142890 892 142896 904
rect 142948 892 142954 944
rect 106182 824 106188 876
rect 106240 864 106246 876
rect 123662 864 123668 876
rect 106240 836 123668 864
rect 106240 824 106246 836
rect 123662 824 123668 836
rect 123720 824 123726 876
rect 123846 824 123852 876
rect 123904 864 123910 876
rect 153102 864 153108 876
rect 123904 836 153108 864
rect 123904 824 123910 836
rect 153102 824 153108 836
rect 153160 824 153166 876
rect 87138 756 87144 808
rect 87196 796 87202 808
rect 110414 796 110420 808
rect 87196 768 110420 796
rect 87196 756 87202 768
rect 110414 756 110420 768
rect 110472 756 110478 808
rect 128354 756 128360 808
rect 128412 796 128418 808
rect 144914 796 144920 808
rect 128412 768 144920 796
rect 128412 756 128418 768
rect 144914 756 144920 768
rect 144972 756 144978 808
rect 84838 688 84844 740
rect 84896 728 84902 740
rect 276014 728 276020 740
rect 84896 700 276020 728
rect 84896 688 84902 700
rect 276014 688 276020 700
rect 276072 688 276078 740
rect 78766 552 78772 604
rect 78824 592 78830 604
rect 237374 592 237380 604
rect 78824 564 237380 592
rect 78824 552 78830 564
rect 237374 552 237380 564
rect 237432 552 237438 604
rect 100754 484 100760 536
rect 100812 524 100818 536
rect 218238 524 218244 536
rect 100812 496 218244 524
rect 100812 484 100818 496
rect 218238 484 218244 496
rect 218296 484 218302 536
rect 117866 416 117872 468
rect 117924 456 117930 468
rect 136266 456 136272 468
rect 117924 428 136272 456
rect 117924 416 117930 428
rect 136266 416 136272 428
rect 136324 416 136330 468
rect 149054 212 149060 264
rect 149112 252 149118 264
rect 256694 252 256700 264
rect 149112 224 256700 252
rect 149112 212 149118 224
rect 256694 212 256700 224
rect 256752 212 256758 264
rect 158714 144 158720 196
rect 158772 184 158778 196
rect 295702 184 295708 196
rect 158772 156 295708 184
rect 158772 144 158778 156
rect 295702 144 295708 156
rect 295760 144 295766 196
rect 79318 76 79324 128
rect 79376 116 79382 128
rect 253658 116 253664 128
rect 79376 88 253664 116
rect 79376 76 79382 88
rect 253658 76 253664 88
rect 253716 76 253722 128
rect 67542 8 67548 60
rect 67600 48 67606 60
rect 126606 48 126612 60
rect 67600 20 126612 48
rect 67600 8 67606 20
rect 126606 8 126612 20
rect 126664 8 126670 60
rect 130286 8 130292 60
rect 130344 48 130350 60
rect 143350 48 143356 60
rect 130344 20 143356 48
rect 130344 8 130350 20
rect 143350 8 143356 20
rect 143408 8 143414 60
rect 178034 8 178040 60
rect 178092 48 178098 60
rect 356514 48 356520 60
rect 178092 20 356520 48
rect 178092 8 178098 20
rect 356514 8 356520 20
rect 356572 8 356578 60
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 89168 700816 89220 700868
rect 96620 700816 96672 700868
rect 95884 700748 95936 700800
rect 154120 700748 154172 700800
rect 24308 700680 24360 700732
rect 100760 700680 100812 700732
rect 8116 700612 8168 700664
rect 99380 700612 99432 700664
rect 87052 700544 87104 700596
rect 283840 700544 283892 700596
rect 84200 700476 84252 700528
rect 348792 700476 348844 700528
rect 80060 700408 80112 700460
rect 413652 700408 413704 700460
rect 77300 700340 77352 700392
rect 478512 700340 478564 700392
rect 74540 700272 74592 700324
rect 543464 700272 543516 700324
rect 72976 699660 73028 699712
rect 76564 699660 76616 699712
rect 217324 699660 217376 699712
rect 218980 699660 219032 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 95240 698912 95292 698964
rect 105452 698912 105504 698964
rect 72424 696940 72476 696992
rect 580172 696940 580224 696992
rect 92572 696192 92624 696244
rect 137836 696192 137888 696244
rect 85580 693404 85632 693456
rect 267648 693404 267700 693456
rect 3424 683204 3476 683256
rect 102140 683204 102192 683256
rect 70492 683136 70544 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 103612 670692 103664 670744
rect 3424 656888 3476 656940
rect 102232 656888 102284 656940
rect 66260 643084 66312 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 104900 632068 104952 632120
rect 67640 630640 67692 630692
rect 579988 630640 580040 630692
rect 3148 618264 3200 618316
rect 107660 618264 107712 618316
rect 64972 616836 65024 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 106280 605820 106332 605872
rect 63500 590656 63552 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 107752 579640 107804 579692
rect 63592 576852 63644 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 110420 565836 110472 565888
rect 62120 563048 62172 563100
rect 580172 563048 580224 563100
rect 3424 553392 3476 553444
rect 109132 553392 109184 553444
rect 59452 536800 59504 536852
rect 579896 536800 579948 536852
rect 3424 527144 3476 527196
rect 111800 527144 111852 527196
rect 60740 524424 60792 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 113180 514768 113232 514820
rect 57980 510620 58032 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 113272 500964 113324 501016
rect 40040 496068 40092 496120
rect 98092 496068 98144 496120
rect 88340 494708 88392 494760
rect 234620 494708 234672 494760
rect 56600 484372 56652 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 114652 474716 114704 474768
rect 58072 470568 58124 470620
rect 580172 470568 580224 470620
rect 3240 462340 3292 462392
rect 117320 462340 117372 462392
rect 55220 456764 55272 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 115940 448536 115992 448588
rect 52460 430584 52512 430636
rect 579896 430584 579948 430636
rect 3424 422288 3476 422340
rect 35164 422288 35216 422340
rect 53932 418140 53984 418192
rect 580172 418140 580224 418192
rect 3148 409844 3200 409896
rect 120172 409844 120224 409896
rect 52552 404336 52604 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 94504 397468 94556 397520
rect 49700 378156 49752 378208
rect 580172 378156 580224 378208
rect 3424 371220 3476 371272
rect 121460 371220 121512 371272
rect 51080 364352 51132 364404
rect 579620 364352 579672 364404
rect 3148 357416 3200 357468
rect 124220 357416 124272 357468
rect 48412 351908 48464 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 122840 345040 122892 345092
rect 46940 324300 46992 324352
rect 580172 324300 580224 324352
rect 3424 318792 3476 318844
rect 124312 318792 124364 318844
rect 47032 311856 47084 311908
rect 579988 311856 580040 311908
rect 3240 304988 3292 305040
rect 126980 304988 127032 305040
rect 45560 298120 45612 298172
rect 580172 298120 580224 298172
rect 3424 292544 3476 292596
rect 125692 292544 125744 292596
rect 42892 271872 42944 271924
rect 580172 271872 580224 271924
rect 3056 266364 3108 266416
rect 128360 266364 128412 266416
rect 44180 258068 44232 258120
rect 580172 258068 580224 258120
rect 3424 253920 3476 253972
rect 129740 253920 129792 253972
rect 41420 244264 41472 244316
rect 580172 244264 580224 244316
rect 3424 240116 3476 240168
rect 129832 240116 129884 240168
rect 40040 231820 40092 231872
rect 579804 231820 579856 231872
rect 41512 218016 41564 218068
rect 579896 218016 579948 218068
rect 3148 213936 3200 213988
rect 131212 213936 131264 213988
rect 38660 205640 38712 205692
rect 580172 205640 580224 205692
rect 3424 201492 3476 201544
rect 133880 201492 133932 201544
rect 35900 191836 35952 191888
rect 580172 191836 580224 191888
rect 3424 187688 3476 187740
rect 132500 187688 132552 187740
rect 37372 178032 37424 178084
rect 580172 178032 580224 178084
rect 91100 173136 91152 173188
rect 217324 173136 217376 173188
rect 89720 171776 89772 171828
rect 201500 171776 201552 171828
rect 76564 170348 76616 170400
rect 96712 170348 96764 170400
rect 83188 168988 83240 169040
rect 331220 168988 331272 169040
rect 80152 167628 80204 167680
rect 396724 167628 396776 167680
rect 35992 165588 36044 165640
rect 580172 165588 580224 165640
rect 76564 164840 76616 164892
rect 462320 164840 462372 164892
rect 3424 162868 3476 162920
rect 135260 162868 135312 162920
rect 33784 162324 33836 162376
rect 119528 162324 119580 162376
rect 20628 162256 20680 162308
rect 151820 162256 151872 162308
rect 2872 162188 2924 162240
rect 153844 162188 153896 162240
rect 1216 162120 1268 162172
rect 188344 162120 188396 162172
rect 3332 162052 3384 162104
rect 196624 162052 196676 162104
rect 17040 161984 17092 162036
rect 220084 161984 220136 162036
rect 12716 161916 12768 161968
rect 233884 161916 233936 161968
rect 4068 161848 4120 161900
rect 285680 161848 285732 161900
rect 8300 161780 8352 161832
rect 302884 161780 302936 161832
rect 8392 161712 8444 161764
rect 305644 161712 305696 161764
rect 2780 161644 2832 161696
rect 309784 161644 309836 161696
rect 15844 161576 15896 161628
rect 422944 161576 422996 161628
rect 7656 161508 7708 161560
rect 449164 161508 449216 161560
rect 69664 161440 69716 161492
rect 557540 161440 557592 161492
rect 69572 160964 69624 161016
rect 201960 160964 202012 161016
rect 12348 160896 12400 160948
rect 150716 160896 150768 160948
rect 12532 160828 12584 160880
rect 152648 160828 152700 160880
rect 2688 160760 2740 160812
rect 174544 160760 174596 160812
rect 35164 160692 35216 160744
rect 118700 160692 118752 160744
rect 119528 160692 119580 160744
rect 295984 160692 296036 160744
rect 3976 160624 4028 160676
rect 215944 160624 215996 160676
rect 3700 160556 3752 160608
rect 246304 160556 246356 160608
rect 73252 160488 73304 160540
rect 353944 160488 353996 160540
rect 2412 160420 2464 160472
rect 283564 160420 283616 160472
rect 20260 160352 20312 160404
rect 336004 160352 336056 160404
rect 13268 160284 13320 160336
rect 381544 160284 381596 160336
rect 3792 160216 3844 160268
rect 400220 160216 400272 160268
rect 3884 160148 3936 160200
rect 445024 160148 445076 160200
rect 2596 160080 2648 160132
rect 463700 160080 463752 160132
rect 5080 159672 5132 159724
rect 20628 159672 20680 159724
rect 18420 159604 18472 159656
rect 33784 159604 33836 159656
rect 73344 159604 73396 159656
rect 156604 159604 156656 159656
rect 6828 159536 6880 159588
rect 12716 159536 12768 159588
rect 16672 159536 16724 159588
rect 150808 159536 150860 159588
rect 9404 159468 9456 159520
rect 152464 159468 152516 159520
rect 11980 159400 12032 159452
rect 161480 159400 161532 159452
rect 6736 159332 6788 159384
rect 180064 159332 180116 159384
rect 6644 159264 6696 159316
rect 251272 159264 251324 159316
rect 6552 159196 6604 159248
rect 267740 159196 267792 159248
rect 940 159128 992 159180
rect 300124 159128 300176 159180
rect 69664 159060 69716 159112
rect 386420 159060 386472 159112
rect 18788 158992 18840 159044
rect 341524 158992 341576 159044
rect 14280 158924 14332 158976
rect 374000 158924 374052 158976
rect 2320 158856 2372 158908
rect 8300 158856 8352 158908
rect 12624 158856 12676 158908
rect 388444 158856 388496 158908
rect 1032 158788 1084 158840
rect 2872 158788 2924 158840
rect 5448 158788 5500 158840
rect 385684 158788 385736 158840
rect 1308 158720 1360 158772
rect 2780 158720 2832 158772
rect 5356 158720 5408 158772
rect 421564 158720 421616 158772
rect 94504 158244 94556 158296
rect 119712 158244 119764 158296
rect 20352 158176 20404 158228
rect 73252 158176 73304 158228
rect 78588 158176 78640 158228
rect 155868 158176 155920 158228
rect 6184 158108 6236 158160
rect 69572 158108 69624 158160
rect 73160 158108 73212 158160
rect 191104 158108 191156 158160
rect 9680 158040 9732 158092
rect 151912 158040 151964 158092
rect 5172 157972 5224 158024
rect 154028 157972 154080 158024
rect 1124 157904 1176 157956
rect 8392 157904 8444 157956
rect 9312 157904 9364 157956
rect 238024 157904 238076 157956
rect 13728 157836 13780 157888
rect 331220 157836 331272 157888
rect 17408 157768 17460 157820
rect 345664 157768 345716 157820
rect 17868 157700 17920 157752
rect 355324 157700 355376 157752
rect 7840 157632 7892 157684
rect 349160 157632 349212 157684
rect 10048 157564 10100 157616
rect 367744 157564 367796 157616
rect 15016 157496 15068 157548
rect 391204 157496 391256 157548
rect 12992 157428 13044 157480
rect 417424 157428 417476 157480
rect 9496 157360 9548 157412
rect 454684 157360 454736 157412
rect 201960 157292 202012 157344
rect 208492 157292 208544 157344
rect 41420 156884 41472 156936
rect 42432 156884 42484 156936
rect 52460 156884 52512 156936
rect 53472 156884 53524 156936
rect 57980 156884 58032 156936
rect 58992 156884 59044 156936
rect 96620 156884 96672 156936
rect 97632 156884 97684 156936
rect 113180 156884 113232 156936
rect 114192 156884 114244 156936
rect 129740 156884 129792 156936
rect 130752 156884 130804 156936
rect 191104 156884 191156 156936
rect 323584 156884 323636 156936
rect 19248 156816 19300 156868
rect 73160 156816 73212 156868
rect 79508 156816 79560 156868
rect 5264 156748 5316 156800
rect 69664 156748 69716 156800
rect 70308 156748 70360 156800
rect 72424 156748 72476 156800
rect 75828 156748 75880 156800
rect 7932 156680 7984 156732
rect 78588 156680 78640 156732
rect 80060 156680 80112 156732
rect 81072 156680 81124 156732
rect 3608 156612 3660 156664
rect 73344 156612 73396 156664
rect 86132 156816 86184 156868
rect 299480 156816 299532 156868
rect 82728 156748 82780 156800
rect 364340 156748 364392 156800
rect 429200 156680 429252 156732
rect 494060 156612 494112 156664
rect 10968 156544 11020 156596
rect 152740 156544 152792 156596
rect 16488 156476 16540 156528
rect 160100 156476 160152 156528
rect 17776 156408 17828 156460
rect 192484 156408 192536 156460
rect 10784 156340 10836 156392
rect 192576 156340 192628 156392
rect 20168 156272 20220 156324
rect 202144 156272 202196 156324
rect 12900 156204 12952 156256
rect 199384 156204 199436 156256
rect 19064 156136 19116 156188
rect 206376 156136 206428 156188
rect 12440 156068 12492 156120
rect 206284 156068 206336 156120
rect 2504 156000 2556 156052
rect 290556 156000 290608 156052
rect 10232 155932 10284 155984
rect 13268 155932 13320 155984
rect 13360 155932 13412 155984
rect 368480 155932 368532 155984
rect 10324 155864 10376 155916
rect 144000 155864 144052 155916
rect 4804 155796 4856 155848
rect 147312 155796 147364 155848
rect 16396 155728 16448 155780
rect 164240 155728 164292 155780
rect 15936 155660 15988 155712
rect 18788 155660 18840 155712
rect 21364 155660 21416 155712
rect 427084 155660 427136 155712
rect 13268 155592 13320 155644
rect 18052 155592 18104 155644
rect 20904 155592 20956 155644
rect 529940 155592 529992 155644
rect 11888 155524 11940 155576
rect 23480 155524 23532 155576
rect 94964 155524 95016 155576
rect 95884 155524 95936 155576
rect 150440 155524 150492 155576
rect 154120 155524 154172 155576
rect 13452 155456 13504 155508
rect 28816 155456 28868 155508
rect 95608 155456 95660 155508
rect 140780 155456 140832 155508
rect 12256 155388 12308 155440
rect 94320 155388 94372 155440
rect 95700 155388 95752 155440
rect 156512 155388 156564 155440
rect 7748 155320 7800 155372
rect 12624 155320 12676 155372
rect 35256 155320 35308 155372
rect 151176 155320 151228 155372
rect 18328 155252 18380 155304
rect 137376 155252 137428 155304
rect 150532 155252 150584 155304
rect 156696 155252 156748 155304
rect 163504 155252 163556 155304
rect 287704 155252 287756 155304
rect 34152 155184 34204 155236
rect 153108 155184 153160 155236
rect 155868 155184 155920 155236
rect 337384 155184 337436 155236
rect 18512 155116 18564 155168
rect 140964 155116 141016 155168
rect 12072 155048 12124 155100
rect 138020 155048 138072 155100
rect 14372 154980 14424 155032
rect 142896 154980 142948 155032
rect 17224 154912 17276 154964
rect 146300 154912 146352 154964
rect 143356 154844 143408 154896
rect 184940 154844 184992 154896
rect 26240 154776 26292 154828
rect 31024 154776 31076 154828
rect 140872 154776 140924 154828
rect 171140 154776 171192 154828
rect 14648 154708 14700 154760
rect 27528 154708 27580 154760
rect 137192 154708 137244 154760
rect 152924 154708 152976 154760
rect 9588 154640 9640 154692
rect 12992 154640 13044 154692
rect 16304 154640 16356 154692
rect 22192 154640 22244 154692
rect 30196 154640 30248 154692
rect 96528 154640 96580 154692
rect 146760 154640 146812 154692
rect 151452 154640 151504 154692
rect 8116 154572 8168 154624
rect 9680 154572 9732 154624
rect 10876 154572 10928 154624
rect 26240 154572 26292 154624
rect 8300 154504 8352 154556
rect 12348 154504 12400 154556
rect 19616 154504 19668 154556
rect 28908 154572 28960 154624
rect 35900 154572 35952 154624
rect 36912 154572 36964 154624
rect 140780 154572 140832 154624
rect 152832 154640 152884 154692
rect 8944 154232 8996 154284
rect 145104 154232 145156 154284
rect 10416 154164 10468 154216
rect 35716 154164 35768 154216
rect 94320 154164 94372 154216
rect 150532 154164 150584 154216
rect 9220 154096 9272 154148
rect 10048 154096 10100 154148
rect 12164 154096 12216 154148
rect 30288 154096 30340 154148
rect 34428 154096 34480 154148
rect 95700 154096 95752 154148
rect 153108 154096 153160 154148
rect 164792 154096 164844 154148
rect 30932 154028 30984 154080
rect 95148 154028 95200 154080
rect 96528 154028 96580 154080
rect 143448 154028 143500 154080
rect 160100 154028 160152 154080
rect 195612 154028 195664 154080
rect 290556 154028 290608 154080
rect 317420 154028 317472 154080
rect 35808 153960 35860 154012
rect 137284 153960 137336 154012
rect 138020 153960 138072 154012
rect 151360 153960 151412 154012
rect 156604 153960 156656 154012
rect 208400 153960 208452 154012
rect 208492 153960 208544 154012
rect 292488 153960 292540 154012
rect 23480 153892 23532 153944
rect 32956 153892 33008 153944
rect 33048 153892 33100 153944
rect 150440 153892 150492 153944
rect 156512 153892 156564 153944
rect 359464 153892 359516 153944
rect 8208 153824 8260 153876
rect 17868 153824 17920 153876
rect 18144 153824 18196 153876
rect 34152 153824 34204 153876
rect 35624 153824 35676 153876
rect 409144 153824 409196 153876
rect 427084 153824 427136 153876
rect 485044 153824 485096 153876
rect 7564 153756 7616 153808
rect 141792 153756 141844 153808
rect 3240 153688 3292 153740
rect 138480 153688 138532 153740
rect 17684 153620 17736 153672
rect 156604 153620 156656 153672
rect 17500 153552 17552 153604
rect 427084 153552 427136 153604
rect 17592 153484 17644 153536
rect 431224 153484 431276 153536
rect 23204 153416 23256 153468
rect 34980 153416 35032 153468
rect 137100 153416 137152 153468
rect 578884 153416 578936 153468
rect 18788 153348 18840 153400
rect 462964 153348 463016 153400
rect 2228 153280 2280 153332
rect 7656 153280 7708 153332
rect 18696 153280 18748 153332
rect 489920 153280 489972 153332
rect 6460 153212 6512 153264
rect 9404 153212 9456 153264
rect 17868 153212 17920 153264
rect 525800 153212 525852 153264
rect 848 153144 900 153196
rect 3332 153144 3384 153196
rect 15108 153144 15160 153196
rect 15844 153144 15896 153196
rect 17132 153144 17184 153196
rect 20352 153144 20404 153196
rect 27528 153144 27580 153196
rect 30932 153144 30984 153196
rect 31024 153144 31076 153196
rect 35808 153144 35860 153196
rect 19892 153076 19944 153128
rect 28816 153076 28868 153128
rect 33048 153076 33100 153128
rect 140872 153144 140924 153196
rect 30196 153008 30248 153060
rect 16028 152940 16080 152992
rect 20628 152940 20680 152992
rect 30288 152940 30340 152992
rect 35716 153008 35768 153060
rect 137192 153076 137244 153128
rect 137284 153076 137336 153128
rect 146760 153076 146812 153128
rect 16212 152872 16264 152924
rect 21364 152872 21416 152924
rect 32956 152872 33008 152924
rect 95608 153008 95660 153060
rect 14924 152736 14976 152788
rect 20904 152736 20956 152788
rect 143448 152668 143500 152720
rect 152004 152668 152056 152720
rect 164792 152668 164844 152720
rect 175280 152668 175332 152720
rect 8024 152600 8076 152652
rect 17408 152600 17460 152652
rect 150532 152600 150584 152652
rect 166264 152600 166316 152652
rect 4988 152532 5040 152584
rect 16672 152532 16724 152584
rect 150440 152532 150492 152584
rect 178040 152532 178092 152584
rect 4896 152464 4948 152516
rect 12532 152464 12584 152516
rect 15752 152464 15804 152516
rect 34428 152464 34480 152516
rect 35348 152464 35400 152516
rect 150992 152464 151044 152516
rect 156696 152464 156748 152516
rect 323032 152464 323084 152516
rect 359464 152464 359516 152516
rect 406384 152464 406436 152516
rect 485044 152464 485096 152516
rect 516784 152464 516836 152516
rect 18880 152260 18932 152312
rect 467104 152260 467156 152312
rect 12992 152192 13044 152244
rect 139584 152192 139636 152244
rect 3424 152124 3476 152176
rect 136272 152124 136324 152176
rect 18604 152056 18656 152108
rect 363604 152056 363656 152108
rect 11796 151988 11848 152040
rect 18144 151988 18196 152040
rect 18972 151988 19024 152040
rect 453304 151988 453356 152040
rect 11704 151920 11756 151972
rect 18420 151920 18472 151972
rect 19984 151920 20036 151972
rect 458824 151920 458876 151972
rect 10692 151852 10744 151904
rect 19892 151852 19944 151904
rect 20076 151852 20128 151904
rect 460204 151852 460256 151904
rect 13176 151716 13228 151768
rect 18236 151784 18288 151836
rect 317420 151716 317472 151768
rect 327724 151716 327776 151768
rect 292488 151648 292540 151700
rect 319444 151648 319496 151700
rect 323584 151648 323636 151700
rect 377404 151648 377456 151700
rect 150900 151580 150952 151632
rect 182180 151580 182232 151632
rect 206376 151580 206428 151632
rect 324412 151580 324464 151632
rect 337384 151580 337436 151632
rect 403624 151580 403676 151632
rect 152924 151512 152976 151564
rect 193220 151512 193272 151564
rect 195612 151512 195664 151564
rect 338120 151512 338172 151564
rect 152832 151444 152884 151496
rect 207020 151444 207072 151496
rect 208400 151444 208452 151496
rect 292672 151444 292724 151496
rect 323032 151444 323084 151496
rect 476764 151444 476816 151496
rect 151360 151376 151412 151428
rect 189080 151376 189132 151428
rect 192576 151376 192628 151428
rect 356704 151376 356756 151428
rect 152004 151308 152056 151360
rect 202880 151308 202932 151360
rect 206284 151308 206336 151360
rect 394700 151308 394752 151360
rect 152096 151240 152148 151292
rect 200120 151240 200172 151292
rect 202144 151240 202196 151292
rect 399484 151240 399536 151292
rect 422944 151240 422996 151292
rect 435364 151240 435416 151292
rect 151452 151172 151504 151224
rect 195980 151172 196032 151224
rect 199384 151172 199436 151224
rect 503720 151172 503772 151224
rect 151268 151104 151320 151156
rect 491944 151104 491996 151156
rect 16120 151036 16172 151088
rect 19800 151036 19852 151088
rect 150992 151036 151044 151088
rect 561680 151036 561732 151088
rect 10600 150560 10652 150612
rect 15936 150560 15988 150612
rect 9036 150492 9088 150544
rect 11980 150492 12032 150544
rect 17316 150492 17368 150544
rect 19616 150492 19668 150544
rect 192484 150492 192536 150544
rect 197360 150492 197412 150544
rect 7656 150424 7708 150476
rect 9128 150424 9180 150476
rect 9312 150424 9364 150476
rect 12900 150424 12952 150476
rect 13084 150424 13136 150476
rect 14464 150424 14516 150476
rect 17408 150424 17460 150476
rect 19708 150424 19760 150476
rect 196624 150424 196676 150476
rect 201500 150424 201552 150476
rect 355324 150424 355376 150476
rect 359464 150424 359516 150476
rect 3424 150356 3476 150408
rect 18328 150356 18380 150408
rect 154120 149812 154172 149864
rect 278044 149812 278096 149864
rect 154028 149744 154080 149796
rect 313924 149744 313976 149796
rect 15936 149676 15988 149728
rect 17040 149676 17092 149728
rect 152740 149676 152792 149728
rect 350540 149676 350592 149728
rect 6368 149064 6420 149116
rect 8300 149064 8352 149116
rect 9128 149064 9180 149116
rect 10232 149064 10284 149116
rect 14464 149064 14516 149116
rect 15752 149064 15804 149116
rect 11980 147636 12032 147688
rect 14280 147636 14332 147688
rect 151176 139340 151228 139392
rect 580172 139340 580224 139392
rect 3516 135804 3568 135856
rect 4896 135804 4948 135856
rect 4896 134580 4948 134632
rect 6184 134580 6236 134632
rect 156696 126896 156748 126948
rect 580172 126896 580224 126948
rect 162124 113092 162176 113144
rect 580172 113092 580224 113144
rect 151084 100648 151136 100700
rect 580172 100648 580224 100700
rect 3148 97928 3200 97980
rect 18512 97928 18564 97980
rect 153936 86912 153988 86964
rect 580172 86912 580224 86964
rect 2964 85484 3016 85536
rect 12992 85484 13044 85536
rect 12992 82832 13044 82884
rect 17132 82832 17184 82884
rect 152648 75828 152700 75880
rect 156696 75828 156748 75880
rect 156604 74332 156656 74384
rect 160100 74332 160152 74384
rect 160744 73108 160796 73160
rect 579988 73108 580040 73160
rect 3424 71612 3476 71664
rect 7564 71612 7616 71664
rect 576124 60664 576176 60716
rect 580172 60664 580224 60716
rect 3332 59304 3384 59356
rect 10324 59304 10376 59356
rect 10324 56924 10376 56976
rect 11704 56924 11756 56976
rect 152556 46860 152608 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 14372 45500 14424 45552
rect 278044 41012 278096 41064
rect 282920 41012 282972 41064
rect 283564 39992 283616 40044
rect 287796 39992 287848 40044
rect 287704 38564 287756 38616
rect 295340 38564 295392 38616
rect 295984 36524 296036 36576
rect 300676 36524 300728 36576
rect 282920 36252 282972 36304
rect 287060 36252 287112 36304
rect 287796 35572 287848 35624
rect 295432 35572 295484 35624
rect 300124 35028 300176 35080
rect 303252 35028 303304 35080
rect 302884 33804 302936 33856
rect 305000 33804 305052 33856
rect 295340 33736 295392 33788
rect 299848 33736 299900 33788
rect 157984 33056 158036 33108
rect 580172 33056 580224 33108
rect 3424 32580 3476 32632
rect 8944 32580 8996 32632
rect 300676 32580 300728 32632
rect 302516 32580 302568 32632
rect 152464 32376 152516 32428
rect 165896 32376 165948 32428
rect 305644 32376 305696 32428
rect 309232 32376 309284 32428
rect 287060 31696 287112 31748
rect 295340 31696 295392 31748
rect 303252 31696 303304 31748
rect 305092 31696 305144 31748
rect 166264 31356 166316 31408
rect 168472 31356 168524 31408
rect 153844 31084 153896 31136
rect 179420 31084 179472 31136
rect 156696 31016 156748 31068
rect 216036 31016 216088 31068
rect 309784 31016 309836 31068
rect 328092 31016 328144 31068
rect 165896 30268 165948 30320
rect 172520 30268 172572 30320
rect 215944 30268 215996 30320
rect 218060 30268 218112 30320
rect 233884 30268 233936 30320
rect 236000 30268 236052 30320
rect 238024 30268 238076 30320
rect 240140 30268 240192 30320
rect 385684 30268 385736 30320
rect 388536 30268 388588 30320
rect 327724 29724 327776 29776
rect 341616 29724 341668 29776
rect 305000 29656 305052 29708
rect 327816 29656 327868 29708
rect 180064 29588 180116 29640
rect 193312 29588 193364 29640
rect 246304 29588 246356 29640
rect 253940 29588 253992 29640
rect 295432 29588 295484 29640
rect 354036 29588 354088 29640
rect 220084 28908 220136 28960
rect 222200 28908 222252 28960
rect 328092 28568 328144 28620
rect 336096 28568 336148 28620
rect 299848 28500 299900 28552
rect 349804 28500 349856 28552
rect 353944 28500 353996 28552
rect 381636 28500 381688 28552
rect 305092 28432 305144 28484
rect 359556 28432 359608 28484
rect 302516 28364 302568 28416
rect 377956 28364 378008 28416
rect 295340 28296 295392 28348
rect 371884 28296 371936 28348
rect 388444 28296 388496 28348
rect 400036 28296 400088 28348
rect 309232 28228 309284 28280
rect 395344 28228 395396 28280
rect 406384 27548 406436 27600
rect 409052 27548 409104 27600
rect 17040 27072 17092 27124
rect 17316 27072 17368 27124
rect 17500 26732 17552 26784
rect 17684 26732 17736 26784
rect 153292 26664 153344 26716
rect 255964 26664 256016 26716
rect 157248 26596 157300 26648
rect 291844 26596 291896 26648
rect 152096 26528 152148 26580
rect 318064 26528 318116 26580
rect 159364 26460 159416 26512
rect 345020 26460 345072 26512
rect 157340 26392 157392 26444
rect 355324 26392 355376 26444
rect 156972 26324 157024 26376
rect 509884 26324 509936 26376
rect 154948 26256 155000 26308
rect 510620 26256 510672 26308
rect 409144 26052 409196 26104
rect 413468 26052 413520 26104
rect 341616 25916 341668 25968
rect 346308 25916 346360 25968
rect 371884 25576 371936 25628
rect 380900 25576 380952 25628
rect 345020 25508 345072 25560
rect 485044 25508 485096 25560
rect 160192 25304 160244 25356
rect 303620 25304 303672 25356
rect 153384 25236 153436 25288
rect 328000 25236 328052 25288
rect 156052 25168 156104 25220
rect 355876 25168 355928 25220
rect 156604 25100 156656 25152
rect 403900 25100 403952 25152
rect 152924 25032 152976 25084
rect 445760 25032 445812 25084
rect 157892 24964 157944 25016
rect 488540 24964 488592 25016
rect 159456 24896 159508 24948
rect 494704 24896 494756 24948
rect 153108 24828 153160 24880
rect 556160 24828 556212 24880
rect 388536 24624 388588 24676
rect 391296 24624 391348 24676
rect 188344 24148 188396 24200
rect 190460 24148 190512 24200
rect 381544 24148 381596 24200
rect 388352 24148 388404 24200
rect 303620 24080 303672 24132
rect 549260 24080 549312 24132
rect 159548 23944 159600 23996
rect 215300 23944 215352 23996
rect 158076 23876 158128 23928
rect 254032 23876 254084 23928
rect 155776 23808 155828 23860
rect 305644 23808 305696 23860
rect 152832 23740 152884 23792
rect 309140 23740 309192 23792
rect 403624 23740 403676 23792
rect 406660 23740 406712 23792
rect 152648 23400 152700 23452
rect 553400 23672 553452 23724
rect 156696 23604 156748 23656
rect 563060 23604 563112 23656
rect 157064 23536 157116 23588
rect 571340 23536 571392 23588
rect 155132 23468 155184 23520
rect 575480 23468 575532 23520
rect 341524 23400 341576 23452
rect 345756 23400 345808 23452
rect 399484 23400 399536 23452
rect 403624 23400 403676 23452
rect 462964 23400 463016 23452
rect 466736 23400 466788 23452
rect 336004 23264 336056 23316
rect 341616 23264 341668 23316
rect 453304 23128 453356 23180
rect 458180 23128 458232 23180
rect 359464 22992 359516 23044
rect 363696 22992 363748 23044
rect 409052 22992 409104 23044
rect 417516 22992 417568 23044
rect 421564 22992 421616 23044
rect 426808 22992 426860 23044
rect 345664 22924 345716 22976
rect 356796 22924 356848 22976
rect 371976 22924 372028 22976
rect 378048 22924 378100 22976
rect 150900 22856 150952 22908
rect 152096 22856 152148 22908
rect 255964 22856 256016 22908
rect 334624 22856 334676 22908
rect 346308 22856 346360 22908
rect 371240 22856 371292 22908
rect 377956 22856 378008 22908
rect 388536 22856 388588 22908
rect 391204 22856 391256 22908
rect 408592 22856 408644 22908
rect 417424 22856 417476 22908
rect 430580 22856 430632 22908
rect 216036 22788 216088 22840
rect 218152 22788 218204 22840
rect 328000 22788 328052 22840
rect 480904 22788 480956 22840
rect 215300 22720 215352 22772
rect 471428 22720 471480 22772
rect 151360 22652 151412 22704
rect 176752 22652 176804 22704
rect 157432 22584 157484 22636
rect 241428 22584 241480 22636
rect 154028 22516 154080 22568
rect 284300 22516 284352 22568
rect 154212 22448 154264 22500
rect 327080 22448 327132 22500
rect 153016 22380 153068 22432
rect 345848 22380 345900 22432
rect 156512 22312 156564 22364
rect 399576 22312 399628 22364
rect 413468 22312 413520 22364
rect 421012 22312 421064 22364
rect 154304 22244 154356 22296
rect 438860 22244 438912 22296
rect 153936 22176 153988 22228
rect 567200 22176 567252 22228
rect 150992 22108 151044 22160
rect 153108 22108 153160 22160
rect 158168 22108 158220 22160
rect 574100 22108 574152 22160
rect 241428 21428 241480 21480
rect 288440 21428 288492 21480
rect 355876 21428 355928 21480
rect 370504 21428 370556 21480
rect 155960 21360 156012 21412
rect 157892 21360 157944 21412
rect 284300 21360 284352 21412
rect 424968 21360 425020 21412
rect 155684 21292 155736 21344
rect 157064 21292 157116 21344
rect 158260 21292 158312 21344
rect 160192 21292 160244 21344
rect 153844 21224 153896 21276
rect 215300 21224 215352 21276
rect 154396 21156 154448 21208
rect 241428 21156 241480 21208
rect 155868 21088 155920 21140
rect 260748 21088 260800 21140
rect 151452 21020 151504 21072
rect 300768 21020 300820 21072
rect 152556 20952 152608 21004
rect 319536 20952 319588 21004
rect 152004 20884 152056 20936
rect 155132 20884 155184 20936
rect 155224 20884 155276 20936
rect 157248 20884 157300 20936
rect 154488 20816 154540 20868
rect 413928 20884 413980 20936
rect 154120 20748 154172 20800
rect 507124 20816 507176 20868
rect 15936 20612 15988 20664
rect 18512 20612 18564 20664
rect 19064 20612 19116 20664
rect 19800 20612 19852 20664
rect 151268 20612 151320 20664
rect 153292 20680 153344 20732
rect 534724 20748 534776 20800
rect 152372 20612 152424 20664
rect 157984 20680 158036 20732
rect 552020 20680 552072 20732
rect 406660 20612 406712 20664
rect 413284 20612 413336 20664
rect 466736 20612 466788 20664
rect 471336 20612 471388 20664
rect 13084 20544 13136 20596
rect 17684 20544 17736 20596
rect 153292 20544 153344 20596
rect 154948 20544 155000 20596
rect 12992 20476 13044 20528
rect 17132 20476 17184 20528
rect 151544 20272 151596 20324
rect 152924 20272 152976 20324
rect 155500 20136 155552 20188
rect 156972 20136 157024 20188
rect 380900 20136 380952 20188
rect 399484 20136 399536 20188
rect 400036 20136 400088 20188
rect 407028 20136 407080 20188
rect 430580 20136 430632 20188
rect 435548 20136 435600 20188
rect 439504 20136 439556 20188
rect 453304 20136 453356 20188
rect 458180 20136 458232 20188
rect 467196 20136 467248 20188
rect 13268 20068 13320 20120
rect 19708 20068 19760 20120
rect 153108 20068 153160 20120
rect 156604 20068 156656 20120
rect 327816 20068 327868 20120
rect 336004 20068 336056 20120
rect 371240 20068 371292 20120
rect 377588 20068 377640 20120
rect 378048 20068 378100 20120
rect 403716 20068 403768 20120
rect 413928 20068 413980 20120
rect 495440 20068 495492 20120
rect 3148 20000 3200 20052
rect 4804 20000 4856 20052
rect 11888 20000 11940 20052
rect 19616 20000 19668 20052
rect 152740 20000 152792 20052
rect 157800 20000 157852 20052
rect 300768 20000 300820 20052
rect 499580 20000 499632 20052
rect 6368 19932 6420 19984
rect 19892 19932 19944 19984
rect 151084 19932 151136 19984
rect 155868 19932 155920 19984
rect 215300 19932 215352 19984
rect 222936 19932 222988 19984
rect 241428 19932 241480 19984
rect 542360 19932 542412 19984
rect 3608 19864 3660 19916
rect 17776 19796 17828 19848
rect 10416 19728 10468 19780
rect 35808 19728 35860 19780
rect 17040 19660 17092 19712
rect 23480 19660 23532 19712
rect 66444 19796 66496 19848
rect 70676 19660 70728 19712
rect 81440 19660 81492 19712
rect 95240 19796 95292 19848
rect 95930 19796 95982 19848
rect 100944 19796 100996 19848
rect 102002 19796 102054 19848
rect 119850 19864 119902 19916
rect 109224 19796 109276 19848
rect 110282 19796 110334 19848
rect 111984 19796 112036 19848
rect 112674 19796 112726 19848
rect 114652 19796 114704 19848
rect 115434 19796 115486 19848
rect 127440 19796 127492 19848
rect 127900 19796 127952 19848
rect 150900 19864 150952 19916
rect 152464 19864 152516 19916
rect 153384 19864 153436 19916
rect 156788 19864 156840 19916
rect 178132 19864 178184 19916
rect 150624 19796 150676 19848
rect 152556 19796 152608 19848
rect 153752 19796 153804 19848
rect 156512 19796 156564 19848
rect 156604 19796 156656 19848
rect 211068 19796 211120 19848
rect 151176 19728 151228 19780
rect 153016 19728 153068 19780
rect 155316 19728 155368 19780
rect 104440 19660 104492 19712
rect 111156 19660 111208 19712
rect 117412 19660 117464 19712
rect 149060 19660 149112 19712
rect 152464 19660 152516 19712
rect 152556 19660 152608 19712
rect 157248 19660 157300 19712
rect 157708 19728 157760 19780
rect 237380 19728 237432 19780
rect 247040 19660 247092 19712
rect 16304 19592 16356 19644
rect 21364 19592 21416 19644
rect 82820 19592 82872 19644
rect 121552 19592 121604 19644
rect 122012 19592 122064 19644
rect 126796 19592 126848 19644
rect 128452 19592 128504 19644
rect 142620 19592 142672 19644
rect 150440 19592 150492 19644
rect 154212 19592 154264 19644
rect 155960 19592 156012 19644
rect 270408 19592 270460 19644
rect 102600 19524 102652 19576
rect 131120 19524 131172 19576
rect 152188 19524 152240 19576
rect 266360 19524 266412 19576
rect 103704 19456 103756 19508
rect 148324 19456 148376 19508
rect 154580 19456 154632 19508
rect 157708 19456 157760 19508
rect 157800 19456 157852 19508
rect 460296 19456 460348 19508
rect 87972 19388 88024 19440
rect 99196 19388 99248 19440
rect 112536 19388 112588 19440
rect 437480 19388 437532 19440
rect 63408 19320 63460 19372
rect 94228 19320 94280 19372
rect 96528 19320 96580 19372
rect 102968 19320 103020 19372
rect 104808 19320 104860 19372
rect 17592 19252 17644 19304
rect 81440 19252 81492 19304
rect 118424 19320 118476 19372
rect 121920 19320 121972 19372
rect 122104 19320 122156 19372
rect 124956 19320 125008 19372
rect 127440 19320 127492 19372
rect 513380 19320 513432 19372
rect 18604 19184 18656 19236
rect 23388 19184 23440 19236
rect 60096 19184 60148 19236
rect 115296 19184 115348 19236
rect 153660 19252 153712 19304
rect 156052 19252 156104 19304
rect 222936 19252 222988 19304
rect 226432 19252 226484 19304
rect 377404 19252 377456 19304
rect 381912 19252 381964 19304
rect 150440 19184 150492 19236
rect 154304 19184 154356 19236
rect 154580 19184 154632 19236
rect 12072 19116 12124 19168
rect 69388 19116 69440 19168
rect 75000 19116 75052 19168
rect 119344 19116 119396 19168
rect 121920 19116 121972 19168
rect 124588 19116 124640 19168
rect 128176 19116 128228 19168
rect 149060 19116 149112 19168
rect 62304 19048 62356 19100
rect 18788 18980 18840 19032
rect 84384 18980 84436 19032
rect 121552 19048 121604 19100
rect 129556 19048 129608 19100
rect 131120 19048 131172 19100
rect 151084 19048 151136 19100
rect 247040 19048 247092 19100
rect 260840 19048 260892 19100
rect 266360 19048 266412 19100
rect 276020 19048 276072 19100
rect 122472 18980 122524 19032
rect 124864 18980 124916 19032
rect 128360 18980 128412 19032
rect 128544 18980 128596 19032
rect 147680 18980 147732 19032
rect 149244 18980 149296 19032
rect 151268 18980 151320 19032
rect 254032 18980 254084 19032
rect 280436 18980 280488 19032
rect 19800 18912 19852 18964
rect 86776 18912 86828 18964
rect 87696 18912 87748 18964
rect 101128 18912 101180 18964
rect 111616 18912 111668 18964
rect 152832 18912 152884 18964
rect 237380 18912 237432 18964
rect 267832 18912 267884 18964
rect 6552 18844 6604 18896
rect 15660 18844 15712 18896
rect 16212 18844 16264 18896
rect 19064 18844 19116 18896
rect 61200 18844 61252 18896
rect 135352 18844 135404 18896
rect 151268 18844 151320 18896
rect 155776 18844 155828 18896
rect 178132 18844 178184 18896
rect 283380 18844 283432 18896
rect 336096 18844 336148 18896
rect 381544 18844 381596 18896
rect 388352 18844 388404 18896
rect 439228 18844 439280 18896
rect 11796 18776 11848 18828
rect 67180 18776 67232 18828
rect 73528 18776 73580 18828
rect 215300 18776 215352 18828
rect 260748 18776 260800 18828
rect 388444 18776 388496 18828
rect 403900 18776 403952 18828
rect 470600 18776 470652 18828
rect 5080 18708 5132 18760
rect 15384 18708 15436 18760
rect 17500 18708 17552 18760
rect 64972 18708 65024 18760
rect 80520 18708 80572 18760
rect 248512 18708 248564 18760
rect 270408 18708 270460 18760
rect 408500 18708 408552 18760
rect 408592 18708 408644 18760
rect 417424 18708 417476 18760
rect 4988 18640 5040 18692
rect 15200 18640 15252 18692
rect 16120 18640 16172 18692
rect 35992 18640 36044 18692
rect 36176 18640 36228 18692
rect 73804 18640 73856 18692
rect 82176 18640 82228 18692
rect 270500 18640 270552 18692
rect 299388 18640 299440 18692
rect 560300 18640 560352 18692
rect 2412 18572 2464 18624
rect 13360 18572 13412 18624
rect 17684 18572 17736 18624
rect 18696 18572 18748 18624
rect 17316 18504 17368 18556
rect 76104 18572 76156 18624
rect 77760 18572 77812 18624
rect 210056 18572 210108 18624
rect 211068 18572 211120 18624
rect 502984 18572 503036 18624
rect 18052 18436 18104 18488
rect 19156 18436 19208 18488
rect 35808 18504 35860 18556
rect 69940 18504 69992 18556
rect 129096 18504 129148 18556
rect 146944 18504 146996 18556
rect 149152 18504 149204 18556
rect 151912 18504 151964 18556
rect 33508 18436 33560 18488
rect 66444 18436 66496 18488
rect 85396 18436 85448 18488
rect 100852 18436 100904 18488
rect 101312 18436 101364 18488
rect 104992 18436 105044 18488
rect 105176 18436 105228 18488
rect 150532 18436 150584 18488
rect 154488 18436 154540 18488
rect 31668 18368 31720 18420
rect 41604 18368 41656 18420
rect 41788 18368 41840 18420
rect 42892 18368 42944 18420
rect 43076 18368 43128 18420
rect 84936 18368 84988 18420
rect 157432 18368 157484 18420
rect 10508 18300 10560 18352
rect 68836 18300 68888 18352
rect 70584 18300 70636 18352
rect 71228 18300 71280 18352
rect 79968 18300 80020 18352
rect 116676 18300 116728 18352
rect 120080 18300 120132 18352
rect 120724 18300 120776 18352
rect 123116 18300 123168 18352
rect 128452 18300 128504 18352
rect 149060 18300 149112 18352
rect 321560 18300 321612 18352
rect 16396 18232 16448 18284
rect 65524 18232 65576 18284
rect 98092 18232 98144 18284
rect 99012 18232 99064 18284
rect 100852 18232 100904 18284
rect 101404 18232 101456 18284
rect 102140 18232 102192 18284
rect 113824 18232 113876 18284
rect 121000 18232 121052 18284
rect 128360 18232 128412 18284
rect 153016 18232 153068 18284
rect 239588 18232 239640 18284
rect 7840 18164 7892 18216
rect 63408 18164 63460 18216
rect 95148 18164 95200 18216
rect 187608 18164 187660 18216
rect 14648 18096 14700 18148
rect 17776 18096 17828 18148
rect 43168 18096 43220 18148
rect 43628 18096 43680 18148
rect 85488 18096 85540 18148
rect 112444 18096 112496 18148
rect 116032 18096 116084 18148
rect 124312 18096 124364 18148
rect 147772 18096 147824 18148
rect 150624 18096 150676 18148
rect 150900 18096 150952 18148
rect 152188 18096 152240 18148
rect 154212 18096 154264 18148
rect 155868 18096 155920 18148
rect 158444 18096 158496 18148
rect 263140 18096 263192 18148
rect 14556 18028 14608 18080
rect 16948 18028 17000 18080
rect 43076 18028 43128 18080
rect 43444 18028 43496 18080
rect 85764 18028 85816 18080
rect 87972 18028 88024 18080
rect 14464 17960 14516 18012
rect 16764 17960 16816 18012
rect 10600 17892 10652 17944
rect 13268 17892 13320 17944
rect 19984 17892 20036 17944
rect 23112 17892 23164 17944
rect 40776 17892 40828 17944
rect 42064 17892 42116 17944
rect 45560 17892 45612 17944
rect 47124 17892 47176 17944
rect 48504 17892 48556 17944
rect 50712 17892 50764 17944
rect 52184 17892 52236 17944
rect 52460 17892 52512 17944
rect 60648 17892 60700 17944
rect 63316 17892 63368 17944
rect 9404 17824 9456 17876
rect 13360 17824 13412 17876
rect 13452 17824 13504 17876
rect 67732 17824 67784 17876
rect 6644 17756 6696 17808
rect 3516 17688 3568 17740
rect 9220 17552 9272 17604
rect 12164 17756 12216 17808
rect 66628 17756 66680 17808
rect 12256 17688 12308 17740
rect 66076 17688 66128 17740
rect 67732 17688 67784 17740
rect 80336 17892 80388 17944
rect 81440 17892 81492 17944
rect 86776 17892 86828 17944
rect 90364 17892 90416 17944
rect 94596 17892 94648 17944
rect 96712 17892 96764 17944
rect 97908 17892 97960 17944
rect 98736 17892 98788 17944
rect 100116 17892 100168 17944
rect 82728 17824 82780 17876
rect 102140 17824 102192 17876
rect 89720 17756 89772 17808
rect 91468 17756 91520 17808
rect 92572 17756 92624 17808
rect 93124 17756 93176 17808
rect 244556 18028 244608 18080
rect 108304 17892 108356 17944
rect 107384 17824 107436 17876
rect 109592 17824 109644 17876
rect 110512 17824 110564 17876
rect 111892 17824 111944 17876
rect 113824 17960 113876 18012
rect 120724 17960 120776 18012
rect 121552 17960 121604 18012
rect 124036 17960 124088 18012
rect 136088 17960 136140 18012
rect 146208 17960 146260 18012
rect 118240 17892 118292 17944
rect 121368 17892 121420 17944
rect 123208 17892 123260 17944
rect 126520 17892 126572 17944
rect 137284 17892 137336 17944
rect 151176 17960 151228 18012
rect 151452 17960 151504 18012
rect 151912 17892 151964 17944
rect 152004 17892 152056 17944
rect 160192 17960 160244 18012
rect 424968 17892 425020 17944
rect 431316 17892 431368 17944
rect 442264 17892 442316 17944
rect 445484 17892 445536 17944
rect 471336 17892 471388 17944
rect 474004 17892 474056 17944
rect 116584 17824 116636 17876
rect 117872 17824 117924 17876
rect 121276 17824 121328 17876
rect 143448 17824 143500 17876
rect 149060 17824 149112 17876
rect 471428 17824 471480 17876
rect 475384 17824 475436 17876
rect 88064 17688 88116 17740
rect 91560 17688 91612 17740
rect 18236 17620 18288 17672
rect 23480 17620 23532 17672
rect 68284 17620 68336 17672
rect 68376 17620 68428 17672
rect 7656 17484 7708 17536
rect 10692 17484 10744 17536
rect 36176 17552 36228 17604
rect 40040 17552 40092 17604
rect 42708 17552 42760 17604
rect 43352 17552 43404 17604
rect 24860 17484 24912 17536
rect 27712 17484 27764 17536
rect 44456 17484 44508 17536
rect 51264 17552 51316 17604
rect 53104 17552 53156 17604
rect 57520 17552 57572 17604
rect 62028 17552 62080 17604
rect 63960 17552 64012 17604
rect 66076 17552 66128 17604
rect 69296 17552 69348 17604
rect 77024 17620 77076 17672
rect 79416 17620 79468 17672
rect 86592 17620 86644 17672
rect 93124 17620 93176 17672
rect 62948 17484 63000 17536
rect 65524 17484 65576 17536
rect 75184 17484 75236 17536
rect 2228 17416 2280 17468
rect 18144 17416 18196 17468
rect 19340 17416 19392 17468
rect 42984 17416 43036 17468
rect 50344 17416 50396 17468
rect 51816 17416 51868 17468
rect 52736 17416 52788 17468
rect 73896 17416 73948 17468
rect 79140 17552 79192 17604
rect 87512 17552 87564 17604
rect 90088 17552 90140 17604
rect 104256 17756 104308 17808
rect 108396 17756 108448 17808
rect 294604 17756 294656 17808
rect 97908 17688 97960 17740
rect 107752 17688 107804 17740
rect 108948 17688 109000 17740
rect 109132 17688 109184 17740
rect 113088 17688 113140 17740
rect 113732 17688 113784 17740
rect 322756 17756 322808 17808
rect 321560 17688 321612 17740
rect 373264 17688 373316 17740
rect 99472 17620 99524 17672
rect 102324 17620 102376 17672
rect 81992 17484 82044 17536
rect 89260 17484 89312 17536
rect 82176 17416 82228 17468
rect 84292 17416 84344 17468
rect 94136 17552 94188 17604
rect 97080 17552 97132 17604
rect 97264 17552 97316 17604
rect 92848 17484 92900 17536
rect 99288 17484 99340 17536
rect 101128 17552 101180 17604
rect 105360 17552 105412 17604
rect 103060 17484 103112 17536
rect 103428 17484 103480 17536
rect 212816 17620 212868 17672
rect 239588 17620 239640 17672
rect 477408 17620 477460 17672
rect 105728 17552 105780 17604
rect 113364 17552 113416 17604
rect 114008 17552 114060 17604
rect 372620 17552 372672 17604
rect 407028 17552 407080 17604
rect 420920 17552 420972 17604
rect 421012 17552 421064 17604
rect 427636 17552 427688 17604
rect 431224 17552 431276 17604
rect 436008 17552 436060 17604
rect 106832 17484 106884 17536
rect 94136 17416 94188 17468
rect 97540 17416 97592 17468
rect 103612 17416 103664 17468
rect 109684 17416 109736 17468
rect 110144 17416 110196 17468
rect 113732 17416 113784 17468
rect 378048 17484 378100 17536
rect 381636 17484 381688 17536
rect 439412 17484 439464 17536
rect 117688 17416 117740 17468
rect 119528 17416 119580 17468
rect 120448 17416 120500 17468
rect 122288 17416 122340 17468
rect 122380 17416 122432 17468
rect 412640 17416 412692 17468
rect 435364 17416 435416 17468
rect 448704 17416 448756 17468
rect 848 17348 900 17400
rect 13452 17348 13504 17400
rect 15568 17348 15620 17400
rect 42340 17348 42392 17400
rect 45744 17348 45796 17400
rect 65892 17348 65944 17400
rect 66260 17348 66312 17400
rect 71596 17348 71648 17400
rect 75092 17348 75144 17400
rect 80704 17348 80756 17400
rect 81072 17348 81124 17400
rect 87604 17348 87656 17400
rect 90732 17348 90784 17400
rect 97264 17348 97316 17400
rect 97356 17348 97408 17400
rect 111340 17348 111392 17400
rect 113364 17348 113416 17400
rect 422392 17348 422444 17400
rect 426808 17348 426860 17400
rect 454776 17348 454828 17400
rect 9680 17280 9732 17332
rect 41420 17280 41472 17332
rect 43444 17280 43496 17332
rect 44916 17280 44968 17332
rect 47952 17280 48004 17332
rect 50344 17280 50396 17332
rect 54944 17280 54996 17332
rect 61384 17280 61436 17332
rect 61844 17280 61896 17332
rect 99196 17280 99248 17332
rect 100024 17280 100076 17332
rect 109776 17280 109828 17332
rect 112352 17280 112404 17332
rect 438124 17280 438176 17332
rect 36544 17212 36596 17264
rect 45100 17212 45152 17264
rect 48228 17212 48280 17264
rect 52736 17212 52788 17264
rect 2320 17144 2372 17196
rect 8944 17144 8996 17196
rect 9036 17144 9088 17196
rect 20628 17144 20680 17196
rect 25044 17144 25096 17196
rect 43812 17144 43864 17196
rect 47768 17144 47820 17196
rect 49700 17144 49752 17196
rect 49792 17144 49844 17196
rect 60004 17212 60056 17264
rect 60832 17144 60884 17196
rect 103704 17212 103756 17264
rect 104164 17212 104216 17264
rect 111524 17212 111576 17264
rect 118884 17212 118936 17264
rect 65892 17144 65944 17196
rect 72148 17144 72200 17196
rect 78128 17144 78180 17196
rect 82360 17144 82412 17196
rect 88800 17144 88852 17196
rect 91376 17144 91428 17196
rect 95056 17144 95108 17196
rect 101496 17144 101548 17196
rect 10784 17076 10836 17128
rect 26240 17076 26292 17128
rect 42064 17076 42116 17128
rect 46020 17076 46072 17128
rect 48872 17076 48924 17128
rect 54576 17076 54628 17128
rect 56508 17076 56560 17128
rect 65524 17076 65576 17128
rect 65708 17076 65760 17128
rect 73988 17076 74040 17128
rect 88248 17076 88300 17128
rect 93768 17076 93820 17128
rect 95700 17076 95752 17128
rect 114560 17144 114612 17196
rect 120908 17212 120960 17264
rect 471980 17212 472032 17264
rect 126888 17144 126940 17196
rect 104532 17076 104584 17128
rect 114008 17076 114060 17128
rect 121736 17076 121788 17128
rect 142160 17144 142212 17196
rect 143632 17144 143684 17196
rect 151544 17144 151596 17196
rect 160192 17144 160244 17196
rect 233516 17144 233568 17196
rect 476764 17076 476816 17128
rect 480260 17076 480312 17128
rect 7748 17008 7800 17060
rect 18420 17008 18472 17060
rect 42156 17008 42208 17060
rect 45836 17008 45888 17060
rect 48136 17008 48188 17060
rect 50528 17008 50580 17060
rect 53656 17008 53708 17060
rect 54944 17008 54996 17060
rect 71872 17008 71924 17060
rect 95148 17008 95200 17060
rect 102324 17008 102376 17060
rect 108304 17008 108356 17060
rect 110788 17008 110840 17060
rect 117688 17008 117740 17060
rect 126152 17008 126204 17060
rect 131120 17008 131172 17060
rect 146300 17008 146352 17060
rect 149152 17008 149204 17060
rect 417516 17008 417568 17060
rect 423680 17008 423732 17060
rect 438860 17008 438912 17060
rect 441988 17008 442040 17060
rect 6000 16940 6052 16992
rect 40868 16940 40920 16992
rect 44180 16940 44232 16992
rect 46756 16940 46808 16992
rect 48688 16940 48740 16992
rect 54760 16940 54812 16992
rect 64144 16940 64196 16992
rect 82820 16940 82872 16992
rect 83832 16940 83884 16992
rect 84844 16940 84896 16992
rect 91008 16940 91060 16992
rect 97816 16940 97868 16992
rect 100760 16940 100812 16992
rect 112996 16940 113048 16992
rect 114468 16940 114520 16992
rect 122380 16940 122432 16992
rect 17776 16872 17828 16924
rect 72700 16872 72752 16924
rect 73344 16872 73396 16924
rect 85488 16872 85540 16924
rect 91192 16872 91244 16924
rect 93584 16872 93636 16924
rect 93768 16872 93820 16924
rect 106096 16872 106148 16924
rect 113456 16872 113508 16924
rect 120908 16872 120960 16924
rect 20076 16804 20128 16856
rect 27620 16804 27672 16856
rect 43536 16804 43588 16856
rect 45652 16804 45704 16856
rect 51448 16804 51500 16856
rect 56048 16804 56100 16856
rect 67824 16804 67876 16856
rect 70124 16804 70176 16856
rect 85856 16804 85908 16856
rect 91008 16804 91060 16856
rect 91744 16804 91796 16856
rect 96712 16804 96764 16856
rect 97816 16804 97868 16856
rect 101312 16804 101364 16856
rect 102416 16804 102468 16856
rect 106924 16804 106976 16856
rect 115112 16804 115164 16856
rect 117504 16804 117556 16856
rect 437480 16804 437532 16856
rect 441620 16804 441672 16856
rect 43628 16736 43680 16788
rect 46204 16736 46256 16788
rect 52552 16736 52604 16788
rect 55864 16736 55916 16788
rect 66444 16736 66496 16788
rect 67916 16736 67968 16788
rect 81624 16736 81676 16788
rect 84476 16736 84528 16788
rect 111248 16736 111300 16788
rect 242808 16736 242860 16788
rect 39304 16668 39356 16720
rect 45468 16668 45520 16720
rect 61660 16668 61712 16720
rect 66812 16668 66864 16720
rect 71780 16668 71832 16720
rect 940 16600 992 16652
rect 8392 16600 8444 16652
rect 44824 16600 44876 16652
rect 46388 16600 46440 16652
rect 61752 16600 61804 16652
rect 64144 16600 64196 16652
rect 64512 16600 64564 16652
rect 65616 16600 65668 16652
rect 66352 16600 66404 16652
rect 68284 16600 68336 16652
rect 72424 16600 72476 16652
rect 76748 16600 76800 16652
rect 82912 16668 82964 16720
rect 85120 16668 85172 16720
rect 93400 16668 93452 16720
rect 94688 16668 94740 16720
rect 97632 16668 97684 16720
rect 104624 16668 104676 16720
rect 107936 16668 107988 16720
rect 240232 16668 240284 16720
rect 97908 16600 97960 16652
rect 116124 16600 116176 16652
rect 7932 16532 7984 16584
rect 11060 16532 11112 16584
rect 10876 16464 10928 16516
rect 70492 16532 70544 16584
rect 116400 16532 116452 16584
rect 116860 16532 116912 16584
rect 122656 16600 122708 16652
rect 123760 16600 123812 16652
rect 129740 16600 129792 16652
rect 132500 16600 132552 16652
rect 153660 16600 153712 16652
rect 153936 16600 153988 16652
rect 121184 16532 121236 16584
rect 129556 16532 129608 16584
rect 133788 16532 133840 16584
rect 142160 16532 142212 16584
rect 147680 16532 147732 16584
rect 16488 16464 16540 16516
rect 18972 16464 19024 16516
rect 10600 16396 10652 16448
rect 66260 16464 66312 16516
rect 83924 16464 83976 16516
rect 86500 16464 86552 16516
rect 111064 16464 111116 16516
rect 117320 16464 117372 16516
rect 143540 16464 143592 16516
rect 158260 16532 158312 16584
rect 26240 16396 26292 16448
rect 96896 16396 96948 16448
rect 99288 16396 99340 16448
rect 201408 16396 201460 16448
rect 212816 16396 212868 16448
rect 295340 16396 295392 16448
rect 6736 16328 6788 16380
rect 15476 16328 15528 16380
rect 24860 16328 24912 16380
rect 91744 16328 91796 16380
rect 95516 16328 95568 16380
rect 262496 16328 262548 16380
rect 267832 16328 267884 16380
rect 280344 16328 280396 16380
rect 280436 16328 280488 16380
rect 380900 16328 380952 16380
rect 6460 16260 6512 16312
rect 19248 16260 19300 16312
rect 21364 16260 21416 16312
rect 71044 16260 71096 16312
rect 71872 16260 71924 16312
rect 79508 16260 79560 16312
rect 112904 16260 112956 16312
rect 117228 16260 117280 16312
rect 117320 16260 117372 16312
rect 291752 16260 291804 16312
rect 391296 16260 391348 16312
rect 399024 16260 399076 16312
rect 15200 16192 15252 16244
rect 43352 16192 43404 16244
rect 55588 16192 55640 16244
rect 73804 16192 73856 16244
rect 90824 16192 90876 16244
rect 283012 16192 283064 16244
rect 294604 16192 294656 16244
rect 417332 16192 417384 16244
rect 13084 16124 13136 16176
rect 41604 16124 41656 16176
rect 47308 16124 47360 16176
rect 74540 16124 74592 16176
rect 77024 16124 77076 16176
rect 81532 16124 81584 16176
rect 82452 16124 82504 16176
rect 87696 16124 87748 16176
rect 89444 16124 89496 16176
rect 223488 16124 223540 16176
rect 240232 16124 240284 16176
rect 436744 16124 436796 16176
rect 7656 16056 7708 16108
rect 41052 16056 41104 16108
rect 53932 16056 53984 16108
rect 86960 16056 87012 16108
rect 91284 16056 91336 16108
rect 327724 16056 327776 16108
rect 372620 16056 372672 16108
rect 377772 16056 377824 16108
rect 381544 16056 381596 16108
rect 395804 16056 395856 16108
rect 399484 16056 399536 16108
rect 438860 16056 438912 16108
rect 4804 15988 4856 16040
rect 39948 15988 40000 16040
rect 55404 15988 55456 16040
rect 97264 15988 97316 16040
rect 98276 15988 98328 16040
rect 374092 15988 374144 16040
rect 381912 15988 381964 16040
rect 390652 15988 390704 16040
rect 395344 15988 395396 16040
rect 476764 15988 476816 16040
rect 5172 15920 5224 15972
rect 20904 15920 20956 15972
rect 23388 15920 23440 15972
rect 59176 15920 59228 15972
rect 63776 15920 63828 15972
rect 66168 15920 66220 15972
rect 66260 15920 66312 15972
rect 111892 15920 111944 15972
rect 114376 15920 114428 15972
rect 478144 15920 478196 15972
rect 3424 15852 3476 15904
rect 40132 15852 40184 15904
rect 57612 15852 57664 15904
rect 111064 15852 111116 15904
rect 116768 15852 116820 15904
rect 485136 15852 485188 15904
rect 13728 15784 13780 15836
rect 15752 15784 15804 15836
rect 17868 15784 17920 15836
rect 33692 15784 33744 15836
rect 56324 15784 56376 15836
rect 91744 15784 91796 15836
rect 92020 15784 92072 15836
rect 98276 15784 98328 15836
rect 102968 15784 103020 15836
rect 107568 15784 107620 15836
rect 109408 15784 109460 15836
rect 143632 15784 143684 15836
rect 150440 15784 150492 15836
rect 158168 15784 158220 15836
rect 13544 15716 13596 15768
rect 22100 15716 22152 15768
rect 50068 15716 50120 15768
rect 53196 15648 53248 15700
rect 61568 15648 61620 15700
rect 62028 15716 62080 15768
rect 66260 15716 66312 15768
rect 73620 15716 73672 15768
rect 81440 15716 81492 15768
rect 91008 15716 91060 15768
rect 118148 15716 118200 15768
rect 122748 15716 122800 15768
rect 123576 15716 123628 15768
rect 65064 15648 65116 15700
rect 90364 15648 90416 15700
rect 98092 15648 98144 15700
rect 99196 15648 99248 15700
rect 112536 15648 112588 15700
rect 15384 15580 15436 15632
rect 20536 15580 20588 15632
rect 84108 15580 84160 15632
rect 89904 15580 89956 15632
rect 97724 15580 97776 15632
rect 98184 15580 98236 15632
rect 18512 15512 18564 15564
rect 22376 15512 22428 15564
rect 19616 15444 19668 15496
rect 45744 15444 45796 15496
rect 81716 15444 81768 15496
rect 153108 15716 153160 15768
rect 132500 15648 132552 15700
rect 143080 15648 143132 15700
rect 77852 15376 77904 15428
rect 152004 15376 152056 15428
rect 65984 15308 66036 15360
rect 167184 15308 167236 15360
rect 377588 15308 377640 15360
rect 381176 15308 381228 15360
rect 18052 15240 18104 15292
rect 20168 15240 20220 15292
rect 66076 15240 66128 15292
rect 70492 15240 70544 15292
rect 86960 15240 87012 15292
rect 89628 15240 89680 15292
rect 153108 15240 153160 15292
rect 179512 15240 179564 15292
rect 16764 15172 16816 15224
rect 24860 15172 24912 15224
rect 42248 15172 42300 15224
rect 42892 15172 42944 15224
rect 60188 15172 60240 15224
rect 61844 15172 61896 15224
rect 75644 15172 75696 15224
rect 78496 15172 78548 15224
rect 81348 15172 81400 15224
rect 82544 15172 82596 15224
rect 87788 15172 87840 15224
rect 88984 15172 89036 15224
rect 90180 15172 90232 15224
rect 92572 15172 92624 15224
rect 92756 15172 92808 15224
rect 95792 15172 95844 15224
rect 99380 15172 99432 15224
rect 101588 15172 101640 15224
rect 124312 15172 124364 15224
rect 128544 15172 128596 15224
rect 130016 15172 130068 15224
rect 4068 15104 4120 15156
rect 10784 15104 10836 15156
rect 13360 15104 13412 15156
rect 77300 15104 77352 15156
rect 122288 15104 122340 15156
rect 124128 15104 124180 15156
rect 155408 15172 155460 15224
rect 532056 15172 532108 15224
rect 158444 15104 158496 15156
rect 187608 15104 187660 15156
rect 205088 15104 205140 15156
rect 8116 15036 8168 15088
rect 15384 15036 15436 15088
rect 2596 14968 2648 15020
rect 10600 14968 10652 15020
rect 10968 14968 11020 15020
rect 64236 15036 64288 15088
rect 64328 15036 64380 15088
rect 65524 15036 65576 15088
rect 142252 15036 142304 15088
rect 150440 15036 150492 15088
rect 2504 14900 2556 14952
rect 10876 14900 10928 14952
rect 15752 14900 15804 14952
rect 89720 14968 89772 15020
rect 131120 14968 131172 15020
rect 243544 14968 243596 15020
rect 18880 14900 18932 14952
rect 19156 14900 19208 14952
rect 58164 14900 58216 14952
rect 3700 14832 3752 14884
rect 15292 14832 15344 14884
rect 15384 14832 15436 14884
rect 62764 14832 62816 14884
rect 3792 14764 3844 14816
rect 19156 14764 19208 14816
rect 20628 14764 20680 14816
rect 65156 14764 65208 14816
rect 19248 14696 19300 14748
rect 61660 14696 61712 14748
rect 4896 14628 4948 14680
rect 18604 14628 18656 14680
rect 19892 14628 19944 14680
rect 60648 14628 60700 14680
rect 90548 14900 90600 14952
rect 210976 14900 211028 14952
rect 349804 14900 349856 14952
rect 390560 14900 390612 14952
rect 439412 14900 439464 14952
rect 442908 14900 442960 14952
rect 449164 14900 449216 14952
rect 456064 14900 456116 14952
rect 71412 14832 71464 14884
rect 197360 14832 197412 14884
rect 242808 14832 242860 14884
rect 263600 14832 263652 14884
rect 291752 14832 291804 14884
rect 353300 14832 353352 14884
rect 399576 14832 399628 14884
rect 413560 14832 413612 14884
rect 477408 14832 477460 14884
rect 488632 14832 488684 14884
rect 81440 14764 81492 14816
rect 216864 14764 216916 14816
rect 233516 14764 233568 14816
rect 242900 14764 242952 14816
rect 244556 14764 244608 14816
rect 284484 14764 284536 14816
rect 295340 14764 295392 14816
rect 407120 14764 407172 14816
rect 412640 14764 412692 14816
rect 423588 14764 423640 14816
rect 423680 14764 423732 14816
rect 435824 14764 435876 14816
rect 439228 14764 439280 14816
rect 445116 14764 445168 14816
rect 448704 14764 448756 14816
rect 513288 14764 513340 14816
rect 69848 14696 69900 14748
rect 78312 14696 78364 14748
rect 81900 14696 81952 14748
rect 223028 14696 223080 14748
rect 223488 14696 223540 14748
rect 317972 14696 318024 14748
rect 322756 14696 322808 14748
rect 450912 14696 450964 14748
rect 460296 14696 460348 14748
rect 471244 14696 471296 14748
rect 480260 14696 480312 14748
rect 507216 14696 507268 14748
rect 5264 14560 5316 14612
rect 21456 14560 21508 14612
rect 22376 14560 22428 14612
rect 47308 14560 47360 14612
rect 57060 14560 57112 14612
rect 60096 14560 60148 14612
rect 64236 14560 64288 14612
rect 67732 14560 67784 14612
rect 76380 14628 76432 14680
rect 234620 14628 234672 14680
rect 240508 14628 240560 14680
rect 396080 14628 396132 14680
rect 406568 14628 406620 14680
rect 427084 14628 427136 14680
rect 427636 14628 427688 14680
rect 493324 14628 493376 14680
rect 79140 14560 79192 14612
rect 86132 14560 86184 14612
rect 297272 14560 297324 14612
rect 355968 14560 356020 14612
rect 521660 14560 521712 14612
rect 1032 14492 1084 14544
rect 13820 14492 13872 14544
rect 17040 14492 17092 14544
rect 42524 14492 42576 14544
rect 54116 14492 54168 14544
rect 79232 14492 79284 14544
rect 89076 14492 89128 14544
rect 282184 14492 282236 14544
rect 283380 14492 283432 14544
rect 498936 14492 498988 14544
rect 2872 14424 2924 14476
rect 40224 14424 40276 14476
rect 40316 14424 40368 14476
rect 40684 14424 40736 14476
rect 55220 14424 55272 14476
rect 79508 14424 79560 14476
rect 81532 14424 81584 14476
rect 251824 14424 251876 14476
rect 263140 14424 263192 14476
rect 570328 14424 570380 14476
rect 9128 14356 9180 14408
rect 21088 14356 21140 14408
rect 30840 14356 30892 14408
rect 44732 14356 44784 14408
rect 60372 14356 60424 14408
rect 131304 14356 131356 14408
rect 445024 14356 445076 14408
rect 448520 14356 448572 14408
rect 15660 14288 15712 14340
rect 21272 14288 21324 14340
rect 61292 14288 61344 14340
rect 108304 14288 108356 14340
rect 64696 14220 64748 14272
rect 88248 14220 88300 14272
rect 93584 14220 93636 14272
rect 97540 14220 97592 14272
rect 441988 14220 442040 14272
rect 448612 14220 448664 14272
rect 50804 14152 50856 14204
rect 69848 14152 69900 14204
rect 79232 14152 79284 14204
rect 84936 14152 84988 14204
rect 58716 14084 58768 14136
rect 77208 14084 77260 14136
rect 79692 14084 79744 14136
rect 168564 14152 168616 14204
rect 420920 14152 420972 14204
rect 424968 14152 425020 14204
rect 93492 14084 93544 14136
rect 148968 14084 149020 14136
rect 417424 14084 417476 14136
rect 423772 14084 423824 14136
rect 66536 14016 66588 14068
rect 81440 14016 81492 14068
rect 108488 14016 108540 14068
rect 113640 14016 113692 14068
rect 117688 14016 117740 14068
rect 119896 14016 119948 14068
rect 157340 14016 157392 14068
rect 159548 14016 159600 14068
rect 78956 13948 79008 14000
rect 80888 13948 80940 14000
rect 82176 13948 82228 14000
rect 188528 13948 188580 14000
rect 18972 13880 19024 13932
rect 92388 13880 92440 13932
rect 115940 13880 115992 13932
rect 117964 13880 118016 13932
rect 118792 13880 118844 13932
rect 121736 13880 121788 13932
rect 123300 13880 123352 13932
rect 129740 13880 129792 13932
rect 18144 13812 18196 13864
rect 19340 13812 19392 13864
rect 27620 13812 27672 13864
rect 33876 13812 33928 13864
rect 78680 13812 78732 13864
rect 81992 13812 82044 13864
rect 102140 13812 102192 13864
rect 108120 13812 108172 13864
rect 108304 13812 108356 13864
rect 125508 13812 125560 13864
rect 126520 13812 126572 13864
rect 127624 13812 127676 13864
rect 5356 13744 5408 13796
rect 10968 13744 11020 13796
rect 3976 13676 4028 13728
rect 65708 13744 65760 13796
rect 67640 13744 67692 13796
rect 71780 13744 71832 13796
rect 83188 13744 83240 13796
rect 86776 13744 86828 13796
rect 114560 13744 114612 13796
rect 118792 13744 118844 13796
rect 122196 13744 122248 13796
rect 137284 13812 137336 13864
rect 149060 13812 149112 13864
rect 152740 13812 152792 13864
rect 435548 13812 435600 13864
rect 440884 13812 440936 13864
rect 155960 13744 156012 13796
rect 159456 13744 159508 13796
rect 201408 13744 201460 13796
rect 327540 13744 327592 13796
rect 13820 13676 13872 13728
rect 66444 13676 66496 13728
rect 75276 13676 75328 13728
rect 211804 13676 211856 13728
rect 15476 13608 15528 13660
rect 67824 13608 67876 13660
rect 73068 13608 73120 13660
rect 211068 13608 211120 13660
rect 223028 13608 223080 13660
rect 241428 13608 241480 13660
rect 18236 13540 18288 13592
rect 68376 13540 68428 13592
rect 78496 13540 78548 13592
rect 229376 13540 229428 13592
rect 10324 13472 10376 13524
rect 23664 13472 23716 13524
rect 33508 13472 33560 13524
rect 37188 13472 37240 13524
rect 53748 13472 53800 13524
rect 57336 13472 57388 13524
rect 81164 13472 81216 13524
rect 255320 13472 255372 13524
rect 276020 13472 276072 13524
rect 282920 13472 282972 13524
rect 31668 13404 31720 13456
rect 36820 13404 36872 13456
rect 65800 13404 65852 13456
rect 70400 13404 70452 13456
rect 89904 13404 89956 13456
rect 244280 13404 244332 13456
rect 253940 13404 253992 13456
rect 432052 13404 432104 13456
rect 21824 13336 21876 13388
rect 43260 13336 43312 13388
rect 50988 13336 51040 13388
rect 70952 13336 71004 13388
rect 80796 13336 80848 13388
rect 258724 13336 258776 13388
rect 282184 13336 282236 13388
rect 314016 13336 314068 13388
rect 363604 13336 363656 13388
rect 398932 13336 398984 13388
rect 17960 13268 18012 13320
rect 40040 13268 40092 13320
rect 51540 13268 51592 13320
rect 75000 13268 75052 13320
rect 86684 13268 86736 13320
rect 276020 13268 276072 13320
rect 280344 13268 280396 13320
rect 285772 13268 285824 13320
rect 298468 13268 298520 13320
rect 405832 13268 405884 13320
rect 13636 13200 13688 13252
rect 40592 13200 40644 13252
rect 54668 13200 54720 13252
rect 82176 13200 82228 13252
rect 91560 13200 91612 13252
rect 307852 13200 307904 13252
rect 318064 13200 318116 13252
rect 520280 13200 520332 13252
rect 16948 13132 17000 13184
rect 79232 13132 79284 13184
rect 91652 13132 91704 13184
rect 318616 13132 318668 13184
rect 319536 13132 319588 13184
rect 351920 13132 351972 13184
rect 355324 13132 355376 13184
rect 417240 13132 417292 13184
rect 3884 13064 3936 13116
rect 23480 13064 23532 13116
rect 24860 13064 24912 13116
rect 33140 13064 33192 13116
rect 33692 13064 33744 13116
rect 68836 13064 68888 13116
rect 77484 13064 77536 13116
rect 241704 13064 241756 13116
rect 243544 13064 243596 13116
rect 516140 13064 516192 13116
rect 11980 12996 12032 13048
rect 21364 12996 21416 13048
rect 68744 12996 68796 13048
rect 168380 12996 168432 13048
rect 210976 12996 211028 13048
rect 299388 12996 299440 13048
rect 9312 12928 9364 12980
rect 91192 12928 91244 12980
rect 108120 12928 108172 12980
rect 119436 12928 119488 12980
rect 119528 12928 119580 12980
rect 156788 12928 156840 12980
rect 168564 12928 168616 12980
rect 222108 12928 222160 12980
rect 58532 12860 58584 12912
rect 115848 12860 115900 12912
rect 118056 12860 118108 12912
rect 118424 12860 118476 12912
rect 84660 12792 84712 12844
rect 87972 12792 88024 12844
rect 59084 12724 59136 12776
rect 102140 12724 102192 12776
rect 70860 12656 70912 12708
rect 179420 12656 179472 12708
rect 8208 12588 8260 12640
rect 91100 12588 91152 12640
rect 133788 12520 133840 12572
rect 140136 12520 140188 12572
rect 89536 12452 89588 12504
rect 90640 12452 90692 12504
rect 8024 12384 8076 12436
rect 102140 12452 102192 12504
rect 105636 12452 105688 12504
rect 96436 12384 96488 12436
rect 106372 12384 106424 12436
rect 116768 12384 116820 12436
rect 148324 12384 148376 12436
rect 155868 12384 155920 12436
rect 168380 12384 168432 12436
rect 180156 12384 180208 12436
rect 197360 12384 197412 12436
rect 202696 12384 202748 12436
rect 377772 12384 377824 12436
rect 380992 12384 381044 12436
rect 388536 12384 388588 12436
rect 390928 12384 390980 12436
rect 403716 12384 403768 12436
rect 408500 12384 408552 12436
rect 441620 12384 441672 12436
rect 444656 12384 444708 12436
rect 1216 12316 1268 12368
rect 69572 12316 69624 12368
rect 81440 12316 81492 12368
rect 170312 12316 170364 12368
rect 423588 12316 423640 12368
rect 435916 12316 435968 12368
rect 436008 12316 436060 12368
rect 449808 12316 449860 12368
rect 2688 12248 2740 12300
rect 67364 12248 67416 12300
rect 70308 12248 70360 12300
rect 160192 12248 160244 12300
rect 179512 12248 179564 12300
rect 241336 12248 241388 12300
rect 430580 12248 430632 12300
rect 433984 12248 434036 12300
rect 442908 12248 442960 12300
rect 448796 12248 448848 12300
rect 20536 12180 20588 12232
rect 24860 12180 24912 12232
rect 72608 12180 72660 12232
rect 183376 12180 183428 12232
rect 241428 12180 241480 12232
rect 270040 12180 270092 12232
rect 417332 12180 417384 12232
rect 443368 12180 443420 12232
rect 6828 12112 6880 12164
rect 12440 12112 12492 12164
rect 21456 12112 21508 12164
rect 23756 12112 23808 12164
rect 75828 12112 75880 12164
rect 202236 12112 202288 12164
rect 222108 12112 222160 12164
rect 255872 12112 255924 12164
rect 378048 12112 378100 12164
rect 394976 12112 395028 12164
rect 427084 12112 427136 12164
rect 463148 12112 463200 12164
rect 10600 12044 10652 12096
rect 19616 12044 19668 12096
rect 20904 12044 20956 12096
rect 78680 12044 78732 12096
rect 85028 12044 85080 12096
rect 223488 12044 223540 12096
rect 244280 12044 244332 12096
rect 284576 12044 284628 12096
rect 395804 12044 395856 12096
rect 10692 11976 10744 12028
rect 20536 11976 20588 12028
rect 23480 11976 23532 12028
rect 88800 11976 88852 12028
rect 88892 11976 88944 12028
rect 93584 11976 93636 12028
rect 94688 11976 94740 12028
rect 249708 11976 249760 12028
rect 255320 11976 255372 12028
rect 264980 11976 265032 12028
rect 283012 11976 283064 12028
rect 322204 11976 322256 12028
rect 358728 11976 358780 12028
rect 434904 11976 434956 12028
rect 448520 12044 448572 12096
rect 460296 12044 460348 12096
rect 485044 12044 485096 12096
rect 498292 12044 498344 12096
rect 448704 11976 448756 12028
rect 448796 11976 448848 12028
rect 459192 11976 459244 12028
rect 470600 11976 470652 12028
rect 510252 11976 510304 12028
rect 8392 11908 8444 11960
rect 18788 11908 18840 11960
rect 19064 11908 19116 11960
rect 40684 11908 40736 11960
rect 55956 11908 56008 11960
rect 66904 11908 66956 11960
rect 77208 11908 77260 11960
rect 81532 11908 81584 11960
rect 82360 11908 82412 11960
rect 245200 11908 245252 11960
rect 248512 11908 248564 11960
rect 260656 11908 260708 11960
rect 262496 11908 262548 11960
rect 348516 11908 348568 11960
rect 353300 11908 353352 11960
rect 440240 11908 440292 11960
rect 448612 11908 448664 11960
rect 491208 11908 491260 11960
rect 8760 11840 8812 11892
rect 41236 11840 41288 11892
rect 50436 11840 50488 11892
rect 67640 11840 67692 11892
rect 82544 11840 82596 11892
rect 261484 11840 261536 11892
rect 263600 11840 263652 11892
rect 421564 11840 421616 11892
rect 435824 11840 435876 11892
rect 488540 11840 488592 11892
rect 488632 11840 488684 11892
rect 493968 11840 494020 11892
rect 1124 11704 1176 11756
rect 15200 11704 15252 11756
rect 18696 11704 18748 11756
rect 22744 11704 22796 11756
rect 18420 11636 18472 11688
rect 63592 11772 63644 11824
rect 65524 11772 65576 11824
rect 81348 11772 81400 11824
rect 88524 11772 88576 11824
rect 303620 11772 303672 11824
rect 380900 11772 380952 11824
rect 387800 11772 387852 11824
rect 390560 11772 390612 11824
rect 520924 11772 520976 11824
rect 20168 11568 20220 11620
rect 22192 11568 22244 11620
rect 18880 11500 18932 11552
rect 77208 11704 77260 11756
rect 79140 11704 79192 11756
rect 93768 11704 93820 11756
rect 107844 11704 107896 11756
rect 431408 11704 431460 11756
rect 438860 11704 438912 11756
rect 445668 11704 445720 11756
rect 26240 11636 26292 11688
rect 43996 11636 44048 11688
rect 56876 11636 56928 11688
rect 108396 11636 108448 11688
rect 218060 11636 218112 11688
rect 219256 11636 219308 11688
rect 445484 11636 445536 11688
rect 512000 11704 512052 11756
rect 513288 11704 513340 11756
rect 531228 11704 531280 11756
rect 453304 11636 453356 11688
rect 457444 11636 457496 11688
rect 480904 11636 480956 11688
rect 485228 11636 485280 11688
rect 57796 11568 57848 11620
rect 107016 11568 107068 11620
rect 58348 11500 58400 11552
rect 82728 11500 82780 11552
rect 103704 11500 103756 11552
rect 125140 11500 125192 11552
rect 15292 11432 15344 11484
rect 71688 11432 71740 11484
rect 71780 11432 71832 11484
rect 84568 11432 84620 11484
rect 95056 11432 95108 11484
rect 110420 11432 110472 11484
rect 211068 11432 211120 11484
rect 213368 11432 213420 11484
rect 67548 11364 67600 11416
rect 151360 11364 151412 11416
rect 21272 11296 21324 11348
rect 77024 11296 77076 11348
rect 133236 11296 133288 11348
rect 136088 11296 136140 11348
rect 111800 11160 111852 11212
rect 378048 11160 378100 11212
rect 13452 11092 13504 11144
rect 10876 11024 10928 11076
rect 116768 11092 116820 11144
rect 398840 11092 398892 11144
rect 92940 11024 92992 11076
rect 95056 11024 95108 11076
rect 95424 11024 95476 11076
rect 97540 11024 97592 11076
rect 70584 10956 70636 11008
rect 96896 10956 96948 11008
rect 100760 10956 100812 11008
rect 106280 10956 106332 11008
rect 107936 10956 107988 11008
rect 114100 10956 114152 11008
rect 115848 10956 115900 11008
rect 151360 10956 151412 11008
rect 151820 10956 151872 11008
rect 179420 10956 179472 11008
rect 198740 10956 198792 11008
rect 59820 10888 59872 10940
rect 61660 10888 61712 10940
rect 66168 10888 66220 10940
rect 71136 10888 71188 10940
rect 78404 10888 78456 10940
rect 183468 10888 183520 10940
rect 24860 10820 24912 10872
rect 63132 10820 63184 10872
rect 68468 10820 68520 10872
rect 182272 10820 182324 10872
rect 183376 10820 183428 10872
rect 209872 10888 209924 10940
rect 210056 10888 210108 10940
rect 236000 10888 236052 10940
rect 241336 10888 241388 10940
rect 268384 10888 268436 10940
rect 223488 10820 223540 10872
rect 276664 10888 276716 10940
rect 276020 10820 276072 10872
rect 299480 10820 299532 10872
rect 85764 10752 85816 10804
rect 88984 10752 89036 10804
rect 223396 10752 223448 10804
rect 249708 10752 249760 10804
rect 284300 10752 284352 10804
rect 303620 10752 303672 10804
rect 312176 10752 312228 10804
rect 19340 10684 19392 10736
rect 29092 10684 29144 10736
rect 33140 10684 33192 10736
rect 42800 10684 42852 10736
rect 51724 10684 51776 10736
rect 75920 10684 75972 10736
rect 82268 10684 82320 10736
rect 249064 10684 249116 10736
rect 282920 10684 282972 10736
rect 417424 10684 417476 10736
rect 14924 10616 14976 10668
rect 23480 10616 23532 10668
rect 30104 10616 30156 10668
rect 44548 10616 44600 10668
rect 56140 10616 56192 10668
rect 94504 10616 94556 10668
rect 95424 10616 95476 10668
rect 96804 10616 96856 10668
rect 101680 10616 101732 10668
rect 102324 10616 102376 10668
rect 104808 10616 104860 10668
rect 109132 10616 109184 10668
rect 110420 10616 110472 10668
rect 285680 10616 285732 10668
rect 299388 10616 299440 10668
rect 309876 10616 309928 10668
rect 5448 10548 5500 10600
rect 23572 10548 23624 10600
rect 40592 10548 40644 10600
rect 65800 10548 65852 10600
rect 90088 10548 90140 10600
rect 305552 10548 305604 10600
rect 14280 10480 14332 10532
rect 41788 10480 41840 10532
rect 55772 10480 55824 10532
rect 96620 10480 96672 10532
rect 96804 10480 96856 10532
rect 103612 10480 103664 10532
rect 108304 10480 108356 10532
rect 313280 10480 313332 10532
rect 336004 10480 336056 10532
rect 362960 10480 363012 10532
rect 398932 10480 398984 10532
rect 427176 10480 427228 10532
rect 11060 10412 11112 10464
rect 57888 10412 57940 10464
rect 61936 10412 61988 10464
rect 68560 10412 68612 10464
rect 92296 10412 92348 10464
rect 337016 10412 337068 10464
rect 354036 10412 354088 10464
rect 367836 10412 367888 10464
rect 417240 10412 417292 10464
rect 449164 10412 449216 10464
rect 13268 10344 13320 10396
rect 59912 10344 59964 10396
rect 61476 10344 61528 10396
rect 68652 10344 68704 10396
rect 68928 10344 68980 10396
rect 82452 10344 82504 10396
rect 83556 10344 83608 10396
rect 278044 10344 278096 10396
rect 285772 10344 285824 10396
rect 548616 10344 548668 10396
rect 9588 10276 9640 10328
rect 88340 10276 88392 10328
rect 94504 10276 94556 10328
rect 96344 10276 96396 10328
rect 96620 10276 96672 10328
rect 96896 10276 96948 10328
rect 98644 10276 98696 10328
rect 108304 10276 108356 10328
rect 114560 10276 114612 10328
rect 116124 10276 116176 10328
rect 132592 10276 132644 10328
rect 534816 10276 534868 10328
rect 60924 10208 60976 10260
rect 128452 10208 128504 10260
rect 147036 10208 147088 10260
rect 154028 10208 154080 10260
rect 182272 10208 182324 10260
rect 183744 10208 183796 10260
rect 52460 10140 52512 10192
rect 78128 10140 78180 10192
rect 78588 10140 78640 10192
rect 131120 10140 131172 10192
rect 54484 10004 54536 10056
rect 92480 10072 92532 10124
rect 93768 10072 93820 10124
rect 98092 10072 98144 10124
rect 135168 10072 135220 10124
rect 64788 9936 64840 9988
rect 68744 9936 68796 9988
rect 70400 9936 70452 9988
rect 10784 9868 10836 9920
rect 81624 9868 81676 9920
rect 88248 9868 88300 9920
rect 104808 10004 104860 10056
rect 113088 10004 113140 10056
rect 128544 10004 128596 10056
rect 140780 10004 140832 10056
rect 166080 9936 166132 9988
rect 125140 9800 125192 9852
rect 127532 9800 127584 9852
rect 156512 9732 156564 9784
rect 180064 9732 180116 9784
rect 84568 9664 84620 9716
rect 91008 9664 91060 9716
rect 12440 9596 12492 9648
rect 72424 9596 72476 9648
rect 86776 9596 86828 9648
rect 91652 9596 91704 9648
rect 98276 9596 98328 9648
rect 100392 9596 100444 9648
rect 101036 9596 101088 9648
rect 111800 9596 111852 9648
rect 115848 9596 115900 9648
rect 123484 9664 123536 9716
rect 131120 9664 131172 9716
rect 240784 9664 240836 9716
rect 123760 9596 123812 9648
rect 124588 9596 124640 9648
rect 143080 9596 143132 9648
rect 143908 9596 143960 9648
rect 156972 9596 157024 9648
rect 159364 9596 159416 9648
rect 183468 9596 183520 9648
rect 232044 9596 232096 9648
rect 356796 9596 356848 9648
rect 360108 9596 360160 9648
rect 367744 9596 367796 9648
rect 372896 9596 372948 9648
rect 387800 9596 387852 9648
rect 391848 9596 391900 9648
rect 403624 9596 403676 9648
rect 406016 9596 406068 9648
rect 434904 9596 434956 9648
rect 438768 9596 438820 9648
rect 502984 9596 503036 9648
rect 506480 9596 506532 9648
rect 23664 9528 23716 9580
rect 68928 9528 68980 9580
rect 18788 9460 18840 9512
rect 70676 9460 70728 9512
rect 80888 9460 80940 9512
rect 91008 9528 91060 9580
rect 102140 9528 102192 9580
rect 107752 9528 107804 9580
rect 111524 9528 111576 9580
rect 112168 9528 112220 9580
rect 114652 9528 114704 9580
rect 154304 9528 154356 9580
rect 158076 9528 158128 9580
rect 209688 9528 209740 9580
rect 210976 9528 211028 9580
rect 223396 9528 223448 9580
rect 292212 9528 292264 9580
rect 356704 9528 356756 9580
rect 360016 9528 360068 9580
rect 405832 9528 405884 9580
rect 408684 9528 408736 9580
rect 234528 9460 234580 9512
rect 236000 9460 236052 9512
rect 242992 9460 243044 9512
rect 463148 9460 463200 9512
rect 467656 9460 467708 9512
rect 18604 9392 18656 9444
rect 90180 9392 90232 9444
rect 91836 9392 91888 9444
rect 282828 9392 282880 9444
rect 284300 9392 284352 9444
rect 343364 9392 343416 9444
rect 510252 9392 510304 9444
rect 517152 9392 517204 9444
rect 52828 9324 52880 9376
rect 83280 9324 83332 9376
rect 86500 9324 86552 9376
rect 277400 9324 277452 9376
rect 285680 9324 285732 9376
rect 354036 9324 354088 9376
rect 438124 9324 438176 9376
rect 449440 9324 449492 9376
rect 491208 9324 491260 9376
rect 510068 9324 510120 9376
rect 17132 9256 17184 9308
rect 26332 9256 26384 9308
rect 94780 9256 94832 9308
rect 291752 9256 291804 9308
rect 404268 9256 404320 9308
rect 427728 9256 427780 9308
rect 440240 9256 440292 9308
rect 452752 9256 452804 9308
rect 456064 9256 456116 9308
rect 471980 9256 472032 9308
rect 474004 9256 474056 9308
rect 491300 9256 491352 9308
rect 507124 9256 507176 9308
rect 534908 9256 534960 9308
rect 20260 9188 20312 9240
rect 56600 9188 56652 9240
rect 65616 9188 65668 9240
rect 84752 9188 84804 9240
rect 87972 9188 88024 9240
rect 287796 9188 287848 9240
rect 313280 9188 313332 9240
rect 377680 9188 377732 9240
rect 390928 9188 390980 9240
rect 400128 9188 400180 9240
rect 408500 9188 408552 9240
rect 435456 9188 435508 9240
rect 435916 9188 435968 9240
rect 458088 9188 458140 9240
rect 458824 9188 458876 9240
rect 470692 9188 470744 9240
rect 491944 9188 491996 9240
rect 528560 9188 528612 9240
rect 13544 9120 13596 9172
rect 40776 9120 40828 9172
rect 55036 9120 55088 9172
rect 93860 9120 93912 9172
rect 98000 9120 98052 9172
rect 106280 9120 106332 9172
rect 109132 9120 109184 9172
rect 318708 9120 318760 9172
rect 348516 9120 348568 9172
rect 357532 9120 357584 9172
rect 380992 9120 381044 9172
rect 412640 9120 412692 9172
rect 424968 9120 425020 9172
rect 436008 9120 436060 9172
rect 448704 9120 448756 9172
rect 476028 9120 476080 9172
rect 488540 9120 488592 9172
rect 526260 9120 526312 9172
rect 531228 9120 531280 9172
rect 541992 9120 542044 9172
rect 19616 9052 19668 9104
rect 67916 9052 67968 9104
rect 68836 9052 68888 9104
rect 86960 9052 87012 9104
rect 88340 9052 88392 9104
rect 20536 8984 20588 9036
rect 71780 8984 71832 9036
rect 81532 8984 81584 9036
rect 15200 8916 15252 8968
rect 20628 8916 20680 8968
rect 21088 8916 21140 8968
rect 82084 8916 82136 8968
rect 85212 8916 85264 8968
rect 91008 8916 91060 8968
rect 95240 8984 95292 9036
rect 97724 8984 97776 9036
rect 100760 9052 100812 9104
rect 350448 9052 350500 9104
rect 378048 9052 378100 9104
rect 393044 9052 393096 9104
rect 394976 9052 395028 9104
rect 403164 9052 403216 9104
rect 413560 9052 413612 9104
rect 449808 9052 449860 9104
rect 449900 9052 449952 9104
rect 498200 9052 498252 9104
rect 498292 9052 498344 9104
rect 531320 9052 531372 9104
rect 534724 9052 534776 9104
rect 571248 9052 571300 9104
rect 103520 8984 103572 9036
rect 107568 8984 107620 9036
rect 355232 8984 355284 9036
rect 377956 8984 378008 9036
rect 430580 8984 430632 9036
rect 431316 8984 431368 9036
rect 445024 8984 445076 9036
rect 445668 8984 445720 9036
rect 478880 8984 478932 9036
rect 493968 8984 494020 9036
rect 565820 8984 565872 9036
rect 101220 8916 101272 8968
rect 101588 8916 101640 8968
rect 382372 8916 382424 8968
rect 385316 8916 385368 8968
rect 394700 8916 394752 8968
rect 398840 8916 398892 8968
rect 416872 8916 416924 8968
rect 426992 8916 427044 8968
rect 503628 8916 503680 8968
rect 516140 8916 516192 8968
rect 577412 8916 577464 8968
rect 49884 8848 49936 8900
rect 64328 8848 64380 8900
rect 70492 8848 70544 8900
rect 56692 8780 56744 8832
rect 83372 8780 83424 8832
rect 84660 8780 84712 8832
rect 154212 8848 154264 8900
rect 160192 8848 160244 8900
rect 186872 8848 186924 8900
rect 135168 8780 135220 8832
rect 139308 8780 139360 8832
rect 82728 8712 82780 8764
rect 101312 8712 101364 8764
rect 88432 8644 88484 8696
rect 91008 8644 91060 8696
rect 94504 8644 94556 8696
rect 96620 8644 96672 8696
rect 100944 8644 100996 8696
rect 128452 8644 128504 8696
rect 131212 8644 131264 8696
rect 351920 8644 351972 8696
rect 354680 8644 354732 8696
rect 68284 8576 68336 8628
rect 162860 8576 162912 8628
rect 68100 8508 68152 8560
rect 172520 8508 172572 8560
rect 59912 8440 59964 8492
rect 95332 8440 95384 8492
rect 444656 8372 444708 8424
rect 452660 8372 452712 8424
rect 78312 8304 78364 8356
rect 84384 8304 84436 8356
rect 102140 8304 102192 8356
rect 107476 8304 107528 8356
rect 8944 8236 8996 8288
rect 94596 8236 94648 8288
rect 96068 8236 96120 8288
rect 97448 8236 97500 8288
rect 98092 8236 98144 8288
rect 102600 8236 102652 8288
rect 102692 8236 102744 8288
rect 114652 8304 114704 8356
rect 115756 8236 115808 8288
rect 125048 8304 125100 8356
rect 119344 8236 119396 8288
rect 123024 8236 123076 8288
rect 65800 8168 65852 8220
rect 71044 8168 71096 8220
rect 81348 8168 81400 8220
rect 85028 8168 85080 8220
rect 116032 8168 116084 8220
rect 119896 8168 119948 8220
rect 122472 8168 122524 8220
rect 130292 8236 130344 8288
rect 137928 8236 137980 8288
rect 184756 8304 184808 8356
rect 191748 8304 191800 8356
rect 213828 8304 213880 8356
rect 146944 8236 146996 8288
rect 149612 8236 149664 8288
rect 327540 8236 327592 8288
rect 330852 8236 330904 8288
rect 149244 8168 149296 8220
rect 151268 8168 151320 8220
rect 80612 8100 80664 8152
rect 155316 8100 155368 8152
rect 202236 8100 202288 8152
rect 223488 8100 223540 8152
rect 94044 8032 94096 8084
rect 207664 8032 207716 8084
rect 22192 7964 22244 8016
rect 90364 7964 90416 8016
rect 94504 7964 94556 8016
rect 213736 7964 213788 8016
rect 37188 7896 37240 7948
rect 70676 7896 70728 7948
rect 74724 7896 74776 7948
rect 204168 7896 204220 7948
rect 213828 7896 213880 7948
rect 236368 7896 236420 7948
rect 318616 7896 318668 7948
rect 332692 7896 332744 7948
rect 29092 7828 29144 7880
rect 92756 7828 92808 7880
rect 125600 7828 125652 7880
rect 127808 7828 127860 7880
rect 129740 7828 129792 7880
rect 265624 7828 265676 7880
rect 318708 7828 318760 7880
rect 342076 7828 342128 7880
rect 24216 7760 24268 7812
rect 43168 7760 43220 7812
rect 54300 7760 54352 7812
rect 90180 7760 90232 7812
rect 90640 7760 90692 7812
rect 319720 7760 319772 7812
rect 362960 7760 363012 7812
rect 389088 7760 389140 7812
rect 4160 7692 4212 7744
rect 40500 7692 40552 7744
rect 42800 7692 42852 7744
rect 64880 7692 64932 7744
rect 90272 7692 90324 7744
rect 321468 7692 321520 7744
rect 345848 7692 345900 7744
rect 383568 7692 383620 7744
rect 15108 7624 15160 7676
rect 35900 7624 35952 7676
rect 36820 7624 36872 7676
rect 81348 7624 81400 7676
rect 88708 7624 88760 7676
rect 94504 7624 94556 7676
rect 96712 7624 96764 7676
rect 364616 7624 364668 7676
rect 23480 7556 23532 7608
rect 80888 7556 80940 7608
rect 109776 7556 109828 7608
rect 385960 7556 386012 7608
rect 61844 7488 61896 7540
rect 124220 7488 124272 7540
rect 143540 7488 143592 7540
rect 152372 7488 152424 7540
rect 61660 7420 61712 7472
rect 121276 7420 121328 7472
rect 84752 7352 84804 7404
rect 140780 7352 140832 7404
rect 57980 7284 58032 7336
rect 108948 7284 109000 7336
rect 93584 7216 93636 7268
rect 191748 7216 191800 7268
rect 57888 7148 57940 7200
rect 95240 7148 95292 7200
rect 23572 7080 23624 7132
rect 96620 7080 96672 7132
rect 69112 7012 69164 7064
rect 156512 7012 156564 7064
rect 150532 6944 150584 6996
rect 153936 6944 153988 6996
rect 127532 6876 127584 6928
rect 134156 6876 134208 6928
rect 150440 6876 150492 6928
rect 160560 6876 160612 6928
rect 3516 6808 3568 6860
rect 17224 6808 17276 6860
rect 56600 6808 56652 6860
rect 95424 6808 95476 6860
rect 101404 6808 101456 6860
rect 104900 6808 104952 6860
rect 107568 6808 107620 6860
rect 111156 6808 111208 6860
rect 111524 6808 111576 6860
rect 116032 6808 116084 6860
rect 118700 6808 118752 6860
rect 121000 6808 121052 6860
rect 184756 6808 184808 6860
rect 204812 6808 204864 6860
rect 507216 6808 507268 6860
rect 509608 6808 509660 6860
rect 72884 6740 72936 6792
rect 186320 6740 186372 6792
rect 213736 6740 213788 6792
rect 278688 6740 278740 6792
rect 431408 6740 431460 6792
rect 434628 6740 434680 6792
rect 476028 6740 476080 6792
rect 484860 6740 484912 6792
rect 80888 6672 80940 6724
rect 88340 6672 88392 6724
rect 85120 6604 85172 6656
rect 214564 6672 214616 6724
rect 391848 6672 391900 6724
rect 395436 6672 395488 6724
rect 449164 6672 449216 6724
rect 455696 6672 455748 6724
rect 462320 6672 462372 6724
rect 471060 6672 471112 6724
rect 471980 6672 472032 6724
rect 481732 6672 481784 6724
rect 88616 6604 88668 6656
rect 231768 6604 231820 6656
rect 427728 6604 427780 6656
rect 441528 6604 441580 6656
rect 467104 6604 467156 6656
rect 480536 6604 480588 6656
rect 50620 6536 50672 6588
rect 69112 6536 69164 6588
rect 85580 6536 85632 6588
rect 272524 6536 272576 6588
rect 282828 6536 282880 6588
rect 321560 6536 321612 6588
rect 400128 6536 400180 6588
rect 430856 6536 430908 6588
rect 433984 6536 434036 6588
rect 448520 6536 448572 6588
rect 458088 6536 458140 6588
rect 467564 6536 467616 6588
rect 476764 6536 476816 6588
rect 492312 6536 492364 6588
rect 509884 6536 509936 6588
rect 529020 6536 529072 6588
rect 53104 6468 53156 6520
rect 72608 6468 72660 6520
rect 73896 6468 73948 6520
rect 82084 6468 82136 6520
rect 87236 6468 87288 6520
rect 282920 6468 282972 6520
rect 291752 6468 291804 6520
rect 340144 6468 340196 6520
rect 23020 6400 23072 6452
rect 43076 6400 43128 6452
rect 52276 6400 52328 6452
rect 79692 6400 79744 6452
rect 86316 6400 86368 6452
rect 294972 6400 295024 6452
rect 359556 6400 359608 6452
rect 390652 6400 390704 6452
rect 17684 6332 17736 6384
rect 40316 6332 40368 6384
rect 53380 6332 53432 6384
rect 86868 6332 86920 6384
rect 92204 6332 92256 6384
rect 1308 6264 1360 6316
rect 33140 6264 33192 6316
rect 57244 6264 57296 6316
rect 92388 6264 92440 6316
rect 26332 6196 26384 6248
rect 86960 6196 87012 6248
rect 92572 6332 92624 6384
rect 300768 6332 300820 6384
rect 341616 6332 341668 6384
rect 363052 6332 363104 6384
rect 373264 6332 373316 6384
rect 413100 6468 413152 6520
rect 417424 6468 417476 6520
rect 448612 6468 448664 6520
rect 449440 6468 449492 6520
rect 465172 6468 465224 6520
rect 467196 6468 467248 6520
rect 484400 6468 484452 6520
rect 485136 6468 485188 6520
rect 493508 6468 493560 6520
rect 528560 6468 528612 6520
rect 547880 6468 547932 6520
rect 408684 6400 408736 6452
rect 417884 6400 417936 6452
rect 421564 6400 421616 6452
rect 458088 6400 458140 6452
rect 460204 6400 460256 6452
rect 473820 6400 473872 6452
rect 475384 6400 475436 6452
rect 502984 6400 503036 6452
rect 520924 6400 520976 6452
rect 546684 6400 546736 6452
rect 310428 6264 310480 6316
rect 319444 6264 319496 6316
rect 331312 6264 331364 6316
rect 353024 6264 353076 6316
rect 403532 6332 403584 6384
rect 416872 6332 416924 6384
rect 426900 6332 426952 6384
rect 427176 6332 427228 6384
rect 462504 6332 462556 6384
rect 467656 6332 467708 6384
rect 492036 6332 492088 6384
rect 493324 6332 493376 6384
rect 525800 6332 525852 6384
rect 526260 6332 526312 6384
rect 565636 6332 565688 6384
rect 403164 6264 403216 6316
rect 427728 6264 427780 6316
rect 435456 6264 435508 6316
rect 471888 6264 471940 6316
rect 478880 6264 478932 6316
rect 543740 6264 543792 6316
rect 97448 6196 97500 6248
rect 361120 6196 361172 6248
rect 363696 6196 363748 6248
rect 368388 6196 368440 6248
rect 370504 6196 370556 6248
rect 403624 6196 403676 6248
rect 403716 6196 403768 6248
rect 466460 6196 466512 6248
rect 470692 6196 470744 6248
rect 481548 6196 481600 6248
rect 485228 6196 485280 6248
rect 566832 6196 566884 6248
rect 20628 6128 20680 6180
rect 59268 6128 59320 6180
rect 68744 6128 68796 6180
rect 80612 6128 80664 6180
rect 87696 6128 87748 6180
rect 262864 6128 262916 6180
rect 265624 6128 265676 6180
rect 536104 6128 536156 6180
rect 65340 6060 65392 6112
rect 150440 6060 150492 6112
rect 186872 6060 186924 6112
rect 191748 6060 191800 6112
rect 204168 6060 204220 6112
rect 221648 6060 221700 6112
rect 345756 6060 345808 6112
rect 351920 6060 351972 6112
rect 360016 6060 360068 6112
rect 362960 6060 363012 6112
rect 62396 5992 62448 6044
rect 144644 5992 144696 6044
rect 145012 5992 145064 6044
rect 155408 5992 155460 6044
rect 80060 5924 80112 5976
rect 88616 5924 88668 5976
rect 89996 5924 90048 5976
rect 92572 5924 92624 5976
rect 127624 5924 127676 5976
rect 140688 5924 140740 5976
rect 94504 5856 94556 5908
rect 98000 5856 98052 5908
rect 140136 5856 140188 5908
rect 146668 5856 146720 5908
rect 66996 5788 67048 5840
rect 174268 5788 174320 5840
rect 367836 5652 367888 5704
rect 370964 5652 371016 5704
rect 59636 5516 59688 5568
rect 67548 5516 67600 5568
rect 83188 5448 83240 5500
rect 86684 5448 86736 5500
rect 86960 5448 87012 5500
rect 97356 5448 97408 5500
rect 103520 5448 103572 5500
rect 109224 5448 109276 5500
rect 113272 5448 113324 5500
rect 116400 5448 116452 5500
rect 144736 5448 144788 5500
rect 151084 5584 151136 5636
rect 454776 5584 454828 5636
rect 459560 5584 459612 5636
rect 150440 5516 150492 5568
rect 154304 5516 154356 5568
rect 277400 5516 277452 5568
rect 283104 5516 283156 5568
rect 314016 5516 314068 5568
rect 316224 5516 316276 5568
rect 394700 5516 394752 5568
rect 400128 5516 400180 5568
rect 412640 5516 412692 5568
rect 415492 5516 415544 5568
rect 454684 5516 454736 5568
rect 462780 5516 462832 5568
rect 471244 5516 471296 5568
rect 476948 5516 477000 5568
rect 491300 5516 491352 5568
rect 494704 5516 494756 5568
rect 534816 5516 534868 5568
rect 539600 5516 539652 5568
rect 149152 5448 149204 5500
rect 155224 5448 155276 5500
rect 180156 5448 180208 5500
rect 185032 5448 185084 5500
rect 84384 5380 84436 5432
rect 179420 5380 179472 5432
rect 71964 5312 72016 5364
rect 198832 5312 198884 5364
rect 232044 5312 232096 5364
rect 247592 5312 247644 5364
rect 59452 5244 59504 5296
rect 60924 5244 60976 5296
rect 79416 5244 79468 5296
rect 213000 5244 213052 5296
rect 214564 5244 214616 5296
rect 236000 5244 236052 5296
rect 74172 5176 74224 5228
rect 205640 5176 205692 5228
rect 207664 5176 207716 5228
rect 346952 5176 347004 5228
rect 51816 5108 51868 5160
rect 66720 5108 66772 5160
rect 83004 5108 83056 5160
rect 224960 5108 225012 5160
rect 236368 5108 236420 5160
rect 315028 5108 315080 5160
rect 55864 5040 55916 5092
rect 80888 5040 80940 5092
rect 84660 5040 84712 5092
rect 274640 5040 274692 5092
rect 51908 4972 51960 5024
rect 77392 4972 77444 5024
rect 88524 4972 88576 5024
rect 291752 4972 291804 5024
rect 27712 4904 27764 4956
rect 44364 4904 44416 4956
rect 53012 4904 53064 4956
rect 84476 4904 84528 4956
rect 86776 4904 86828 4956
rect 301964 4904 302016 4956
rect 11152 4836 11204 4888
rect 41696 4836 41748 4888
rect 54944 4836 54996 4888
rect 87972 4836 88024 4888
rect 109684 4836 109736 4888
rect 111800 4836 111852 4888
rect 114468 4836 114520 4888
rect 118056 4836 118108 4888
rect 121184 4836 121236 4888
rect 489920 4836 489972 4888
rect 22744 4768 22796 4820
rect 56508 4768 56560 4820
rect 68560 4768 68612 4820
rect 56048 4700 56100 4752
rect 73804 4700 73856 4752
rect 108396 4768 108448 4820
rect 114100 4768 114152 4820
rect 121460 4768 121512 4820
rect 521568 4768 521620 4820
rect 139400 4700 139452 4752
rect 146576 4700 146628 4752
rect 149152 4700 149204 4752
rect 68652 4632 68704 4684
rect 133788 4632 133840 4684
rect 76196 4564 76248 4616
rect 127624 4564 127676 4616
rect 131120 4564 131172 4616
rect 137928 4564 137980 4616
rect 59268 4496 59320 4548
rect 101680 4496 101732 4548
rect 62580 4428 62632 4480
rect 153752 4360 153804 4412
rect 156604 4360 156656 4412
rect 144828 4224 144880 4276
rect 150532 4224 150584 4276
rect 54576 4088 54628 4140
rect 57244 4088 57296 4140
rect 75184 4088 75236 4140
rect 106924 4088 106976 4140
rect 109500 4088 109552 4140
rect 116676 4088 116728 4140
rect 119436 4088 119488 4140
rect 123484 4088 123536 4140
rect 127624 4088 127676 4140
rect 131120 4088 131172 4140
rect 145932 4088 145984 4140
rect 251824 4088 251876 4140
rect 252468 4088 252520 4140
rect 313924 4088 313976 4140
rect 317328 4088 317380 4140
rect 362960 4088 363012 4140
rect 367008 4088 367060 4140
rect 516784 4088 516836 4140
rect 519544 4088 519596 4140
rect 59176 4020 59228 4072
rect 124680 4020 124732 4072
rect 127808 4020 127860 4072
rect 137652 4020 137704 4072
rect 146944 4020 146996 4072
rect 157984 4020 158036 4072
rect 180064 4020 180116 4072
rect 187332 4020 187384 4072
rect 85028 3952 85080 4004
rect 156604 3952 156656 4004
rect 179420 3952 179472 4004
rect 192024 3952 192076 4004
rect 234528 3952 234580 4004
rect 251180 3952 251232 4004
rect 460296 3952 460348 4004
rect 469864 3952 469916 4004
rect 71136 3884 71188 3936
rect 152924 3884 152976 3936
rect 172520 3884 172572 3936
rect 181444 3884 181496 3936
rect 186320 3884 186372 3936
rect 212172 3884 212224 3936
rect 213000 3884 213052 3936
rect 238116 3884 238168 3936
rect 240784 3884 240836 3936
rect 244188 3884 244240 3936
rect 262864 3884 262916 3936
rect 33600 3816 33652 3868
rect 36544 3816 36596 3868
rect 43076 3816 43128 3868
rect 46572 3816 46624 3868
rect 61568 3816 61620 3868
rect 85672 3816 85724 3868
rect 90180 3816 90232 3868
rect 92756 3816 92808 3868
rect 93860 3816 93912 3868
rect 97448 3816 97500 3868
rect 101220 3816 101272 3868
rect 34796 3748 34848 3800
rect 45284 3748 45336 3800
rect 49516 3748 49568 3800
rect 62028 3748 62080 3800
rect 64144 3748 64196 3800
rect 69664 3748 69716 3800
rect 73896 3748 73948 3800
rect 101036 3748 101088 3800
rect 104256 3816 104308 3868
rect 108396 3816 108448 3868
rect 108580 3816 108632 3868
rect 195980 3816 196032 3868
rect 198832 3816 198884 3868
rect 108212 3748 108264 3800
rect 108488 3748 108540 3800
rect 201684 3748 201736 3800
rect 205640 3816 205692 3868
rect 220452 3816 220504 3868
rect 231768 3816 231820 3868
rect 258264 3816 258316 3868
rect 261484 3816 261536 3868
rect 266544 3816 266596 3868
rect 278688 3884 278740 3936
rect 273628 3816 273680 3868
rect 282920 3816 282972 3868
rect 285128 3816 285180 3868
rect 305644 3884 305696 3936
rect 313832 3884 313884 3936
rect 459560 3884 459612 3936
rect 467472 3884 467524 3936
rect 467564 3884 467616 3936
rect 479340 3884 479392 3936
rect 291384 3816 291436 3868
rect 292212 3816 292264 3868
rect 307944 3816 307996 3868
rect 309876 3816 309928 3868
rect 325608 3816 325660 3868
rect 330852 3816 330904 3868
rect 339868 3816 339920 3868
rect 342076 3816 342128 3868
rect 348056 3816 348108 3868
rect 448520 3816 448572 3868
rect 474556 3816 474608 3868
rect 494796 3816 494848 3868
rect 507676 3816 507728 3868
rect 206192 3748 206244 3800
rect 211804 3748 211856 3800
rect 227536 3748 227588 3800
rect 236000 3748 236052 3800
rect 276112 3748 276164 3800
rect 276664 3748 276716 3800
rect 290188 3748 290240 3800
rect 291752 3748 291804 3800
rect 311440 3748 311492 3800
rect 321560 3748 321612 3800
rect 32404 3544 32456 3596
rect 43444 3680 43496 3732
rect 48964 3680 49016 3732
rect 40684 3612 40736 3664
rect 41880 3544 41932 3596
rect 44824 3544 44876 3596
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 12348 3476 12400 3528
rect 13084 3476 13136 3528
rect 38384 3476 38436 3528
rect 42156 3476 42208 3528
rect 49332 3612 49384 3664
rect 57336 3680 57388 3732
rect 89168 3680 89220 3732
rect 92480 3680 92532 3732
rect 93952 3680 94004 3732
rect 50528 3544 50580 3596
rect 52552 3544 52604 3596
rect 58440 3612 58492 3664
rect 61384 3612 61436 3664
rect 92940 3612 92992 3664
rect 60832 3544 60884 3596
rect 66904 3544 66956 3596
rect 103336 3680 103388 3732
rect 103428 3680 103480 3732
rect 200672 3680 200724 3732
rect 204812 3680 204864 3732
rect 233424 3680 233476 3732
rect 242900 3680 242952 3732
rect 244096 3680 244148 3732
rect 244188 3680 244240 3732
rect 248788 3680 248840 3732
rect 249064 3680 249116 3732
rect 272432 3680 272484 3732
rect 272524 3680 272576 3732
rect 293684 3680 293736 3732
rect 300768 3680 300820 3732
rect 322112 3680 322164 3732
rect 327724 3680 327776 3732
rect 330392 3680 330444 3732
rect 331312 3748 331364 3800
rect 342168 3748 342220 3800
rect 452660 3748 452712 3800
rect 466276 3748 466328 3800
rect 466460 3748 466512 3800
rect 497096 3748 497148 3800
rect 333888 3680 333940 3732
rect 334624 3680 334676 3732
rect 344560 3680 344612 3732
rect 96344 3612 96396 3664
rect 104532 3612 104584 3664
rect 107016 3612 107068 3664
rect 115204 3612 115256 3664
rect 116676 3612 116728 3664
rect 214656 3612 214708 3664
rect 224960 3612 225012 3664
rect 277124 3612 277176 3664
rect 284300 3612 284352 3664
rect 285036 3612 285088 3664
rect 285128 3612 285180 3664
rect 304356 3612 304408 3664
rect 310428 3612 310480 3664
rect 336280 3612 336332 3664
rect 340144 3612 340196 3664
rect 352840 3680 352892 3732
rect 370964 3680 371016 3732
rect 379980 3680 380032 3732
rect 389088 3680 389140 3732
rect 394240 3680 394292 3732
rect 430580 3680 430632 3732
rect 434444 3680 434496 3732
rect 448612 3680 448664 3732
rect 514760 3680 514812 3732
rect 351920 3612 351972 3664
rect 359924 3612 359976 3664
rect 377404 3612 377456 3664
rect 388260 3612 388312 3664
rect 388444 3612 388496 3664
rect 402520 3612 402572 3664
rect 403624 3612 403676 3664
rect 420184 3612 420236 3664
rect 438768 3612 438820 3664
rect 460388 3612 460440 3664
rect 462504 3612 462556 3664
rect 533712 3612 533764 3664
rect 96896 3544 96948 3596
rect 102232 3544 102284 3596
rect 102876 3544 102928 3596
rect 103428 3544 103480 3596
rect 105084 3544 105136 3596
rect 108488 3544 108540 3596
rect 108948 3544 109000 3596
rect 81440 3476 81492 3528
rect 88432 3476 88484 3528
rect 108120 3476 108172 3528
rect 108304 3476 108356 3528
rect 109316 3476 109368 3528
rect 111064 3544 111116 3596
rect 114008 3544 114060 3596
rect 117872 3544 117924 3596
rect 433248 3544 433300 3596
rect 436008 3544 436060 3596
rect 440332 3544 440384 3596
rect 440884 3544 440936 3596
rect 452108 3544 452160 3596
rect 452752 3544 452804 3596
rect 456892 3544 456944 3596
rect 457444 3544 457496 3596
rect 537208 3544 537260 3596
rect 543740 3544 543792 3596
rect 551468 3544 551520 3596
rect 116400 3476 116452 3528
rect 118240 3476 118292 3528
rect 468668 3476 468720 3528
rect 473820 3476 473872 3528
rect 501788 3476 501840 3528
rect 503628 3476 503680 3528
rect 505376 3476 505428 3528
rect 509608 3476 509660 3528
rect 523040 3476 523092 3528
rect 525800 3476 525852 3528
rect 554964 3476 555016 3528
rect 562324 3476 562376 3528
rect 564440 3476 564492 3528
rect 571248 3476 571300 3528
rect 573916 3476 573968 3528
rect 5264 3408 5316 3460
rect 17684 3408 17736 3460
rect 20628 3408 20680 3460
rect 40684 3408 40736 3460
rect 43628 3408 43680 3460
rect 45468 3408 45520 3460
rect 47032 3408 47084 3460
rect 47492 3408 47544 3460
rect 48964 3408 49016 3460
rect 50344 3408 50396 3460
rect 51356 3408 51408 3460
rect 54760 3408 54812 3460
rect 56048 3408 56100 3460
rect 60096 3408 60148 3460
rect 110512 3408 110564 3460
rect 113916 3408 113968 3460
rect 475752 3408 475804 3460
rect 492036 3408 492088 3460
rect 581000 3408 581052 3460
rect 42248 3340 42300 3392
rect 50712 3340 50764 3392
rect 54944 3340 54996 3392
rect 35992 3272 36044 3324
rect 39304 3272 39356 3324
rect 49148 3272 49200 3324
rect 59636 3340 59688 3392
rect 79508 3340 79560 3392
rect 98644 3340 98696 3392
rect 84936 3272 84988 3324
rect 91560 3272 91612 3324
rect 92940 3272 92992 3324
rect 96252 3272 96304 3324
rect 97264 3272 97316 3324
rect 99840 3340 99892 3392
rect 60004 3204 60056 3256
rect 63224 3204 63276 3256
rect 82176 3204 82228 3256
rect 95148 3204 95200 3256
rect 98000 3204 98052 3256
rect 104808 3340 104860 3392
rect 108212 3340 108264 3392
rect 121092 3340 121144 3392
rect 121276 3340 121328 3392
rect 128176 3340 128228 3392
rect 131212 3340 131264 3392
rect 135260 3340 135312 3392
rect 149520 3340 149572 3392
rect 151360 3340 151412 3392
rect 39580 3136 39632 3188
rect 42064 3136 42116 3188
rect 92388 3136 92440 3188
rect 111616 3272 111668 3324
rect 111800 3272 111852 3324
rect 117872 3272 117924 3324
rect 146668 3272 146720 3324
rect 155408 3340 155460 3392
rect 160100 3340 160152 3392
rect 161296 3340 161348 3392
rect 174544 3340 174596 3392
rect 176660 3340 176712 3392
rect 184940 3340 184992 3392
rect 186136 3340 186188 3392
rect 299480 3340 299532 3392
rect 300768 3340 300820 3392
rect 307852 3340 307904 3392
rect 309048 3340 309100 3392
rect 354680 3340 354732 3392
rect 358728 3340 358780 3392
rect 358820 3340 358872 3392
rect 362316 3340 362368 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 160560 3272 160612 3324
rect 163688 3272 163740 3324
rect 223488 3272 223540 3324
rect 231032 3272 231084 3324
rect 252468 3272 252520 3324
rect 259460 3272 259512 3324
rect 321468 3272 321520 3324
rect 323308 3272 323360 3324
rect 372620 3272 372672 3324
rect 376484 3272 376536 3324
rect 484400 3272 484452 3324
rect 487620 3272 487672 3324
rect 565820 3272 565872 3324
rect 569132 3272 569184 3324
rect 101312 3204 101364 3256
rect 118792 3204 118844 3256
rect 471888 3204 471940 3256
rect 473452 3204 473504 3256
rect 102600 3136 102652 3188
rect 117596 3136 117648 3188
rect 124588 3136 124640 3188
rect 156972 3136 157024 3188
rect 162860 3136 162912 3188
rect 169576 3136 169628 3188
rect 221648 3136 221700 3188
rect 223948 3136 224000 3188
rect 360108 3136 360160 3188
rect 363512 3136 363564 3188
rect 413284 3136 413336 3188
rect 416688 3136 416740 3188
rect 434628 3136 434680 3188
rect 437940 3136 437992 3188
rect 481548 3136 481600 3188
rect 484032 3136 484084 3188
rect 512644 3136 512696 3188
rect 515956 3136 516008 3188
rect 91744 3068 91796 3120
rect 105728 3068 105780 3120
rect 191748 3068 191800 3120
rect 195612 3068 195664 3120
rect 220728 3068 220780 3120
rect 246396 3068 246448 3120
rect 291844 3068 291896 3120
rect 294880 3068 294932 3120
rect 294972 3068 295024 3120
rect 298468 3068 298520 3120
rect 445116 3068 445168 3120
rect 448612 3068 448664 3120
rect 103980 3000 104032 3052
rect 108580 3000 108632 3052
rect 150440 3000 150492 3052
rect 153844 3000 153896 3052
rect 157340 3000 157392 3052
rect 232228 3000 232280 3052
rect 278044 3000 278096 3052
rect 280712 3000 280764 3052
rect 395436 3000 395488 3052
rect 397736 3000 397788 3052
rect 1676 2932 1728 2984
rect 3424 2932 3476 2984
rect 37188 2932 37240 2984
rect 43536 2932 43588 2984
rect 133788 2932 133840 2984
rect 138848 2932 138900 2984
rect 139400 2932 139452 2984
rect 142436 2932 142488 2984
rect 194968 2932 195020 2984
rect 214472 2932 214524 2984
rect 214564 2932 214616 2984
rect 235816 2932 235868 2984
rect 322204 2932 322256 2984
rect 326804 2932 326856 2984
rect 118608 2864 118660 2916
rect 122288 2864 122340 2916
rect 129740 2864 129792 2916
rect 141240 2864 141292 2916
rect 154488 2864 154540 2916
rect 157800 2864 157852 2916
rect 201040 2864 201092 2916
rect 221556 2864 221608 2916
rect 258724 2864 258776 2916
rect 262956 2864 263008 2916
rect 363052 2864 363104 2916
rect 365812 2864 365864 2916
rect 368388 2864 368440 2916
rect 370596 2864 370648 2916
rect 115848 2796 115900 2848
rect 33140 2728 33192 2780
rect 112168 2728 112220 2780
rect 112444 2728 112496 2780
rect 114468 2728 114520 2780
rect 144736 2796 144788 2848
rect 153016 2796 153068 2848
rect 158904 2796 158956 2848
rect 202788 2796 202840 2848
rect 208584 2796 208636 2848
rect 218152 2796 218204 2848
rect 225144 2796 225196 2848
rect 247040 2796 247092 2848
rect 249984 2796 250036 2848
rect 274640 2796 274692 2848
rect 279516 2796 279568 2848
rect 409788 2796 409840 2848
rect 411904 2796 411956 2848
rect 427728 2796 427780 2848
rect 429660 2796 429712 2848
rect 445668 2796 445720 2848
rect 447416 2796 447468 2848
rect 521568 2796 521620 2848
rect 524236 2796 524288 2848
rect 552572 2796 552624 2848
rect 559748 2796 559800 2848
rect 149612 2728 149664 2780
rect 572720 2796 572772 2848
rect 76564 2660 76616 2712
rect 214564 2660 214616 2712
rect 214656 2660 214708 2712
rect 445668 2660 445720 2712
rect 116584 2592 116636 2644
rect 117872 2592 117924 2644
rect 124220 2592 124272 2644
rect 130568 2592 130620 2644
rect 143908 2592 143960 2644
rect 153752 2592 153804 2644
rect 195980 2592 196032 2644
rect 409788 2592 409840 2644
rect 78220 2524 78272 2576
rect 220728 2524 220780 2576
rect 58900 2456 58952 2508
rect 118608 2456 118660 2508
rect 76012 2388 76064 2440
rect 157340 2456 157392 2508
rect 173532 2456 173584 2508
rect 202788 2456 202840 2508
rect 158812 2388 158864 2440
rect 218152 2388 218204 2440
rect 237380 2388 237432 2440
rect 247040 2388 247092 2440
rect 67916 2320 67968 2372
rect 112076 2320 112128 2372
rect 120724 2320 120776 2372
rect 274824 2320 274876 2372
rect 87604 2252 87656 2304
rect 264152 2252 264204 2304
rect 81440 2184 81492 2236
rect 87144 2184 87196 2236
rect 91652 2184 91704 2236
rect 278320 2184 278372 2236
rect 60740 2116 60792 2168
rect 132960 2116 133012 2168
rect 135076 2116 135128 2168
rect 144828 2116 144880 2168
rect 144920 2116 144972 2168
rect 194968 2116 195020 2168
rect 200672 2116 200724 2168
rect 404820 2116 404872 2168
rect 63500 2048 63552 2100
rect 74356 1980 74408 2032
rect 106188 1980 106240 2032
rect 112536 1980 112588 2032
rect 129740 1980 129792 2032
rect 75460 1912 75512 1964
rect 100760 1912 100812 1964
rect 104808 1912 104860 1964
rect 121460 1912 121512 1964
rect 153108 2048 153160 2100
rect 201040 2048 201092 2100
rect 201684 2048 201736 2100
rect 418988 2048 419040 2100
rect 140780 1980 140832 2032
rect 154488 1980 154540 2032
rect 151820 1912 151872 1964
rect 97540 1844 97592 1896
rect 115848 1844 115900 1896
rect 80704 1776 80756 1828
rect 150440 1776 150492 1828
rect 121184 1640 121236 1692
rect 124128 1640 124180 1692
rect 137284 1640 137336 1692
rect 178040 1640 178092 1692
rect 121368 1572 121420 1624
rect 128360 1572 128412 1624
rect 122840 1504 122892 1556
rect 124864 1504 124916 1556
rect 122748 1436 122800 1488
rect 125876 1436 125928 1488
rect 142804 1572 142856 1624
rect 136548 1504 136600 1556
rect 146300 1504 146352 1556
rect 85948 1232 86000 1284
rect 122932 1368 122984 1420
rect 123024 1368 123076 1420
rect 133788 1436 133840 1488
rect 140044 1436 140096 1488
rect 115848 1300 115900 1352
rect 121184 1300 121236 1352
rect 126980 1300 127032 1352
rect 136272 1368 136324 1420
rect 149060 1436 149112 1488
rect 218244 1436 218296 1488
rect 228732 1436 228784 1488
rect 142896 1368 142948 1420
rect 137284 1300 137336 1352
rect 158720 1368 158772 1420
rect 148324 1300 148376 1352
rect 150808 1300 150860 1352
rect 114468 1232 114520 1284
rect 121368 1232 121420 1284
rect 121460 1232 121512 1284
rect 129648 1232 129700 1284
rect 146300 1232 146352 1284
rect 149244 1232 149296 1284
rect 64880 1164 64932 1216
rect 114100 1164 114152 1216
rect 139492 1164 139544 1216
rect 153016 1164 153068 1216
rect 77116 1096 77168 1148
rect 239312 1368 239364 1420
rect 276020 1368 276072 1420
rect 281908 1368 281960 1420
rect 313280 1368 313332 1420
rect 320916 1368 320968 1420
rect 72332 1028 72384 1080
rect 173532 1028 173584 1080
rect 69664 960 69716 1012
rect 133788 960 133840 1012
rect 142804 960 142856 1012
rect 158812 960 158864 1012
rect 60924 892 60976 944
rect 122748 892 122800 944
rect 122932 892 122984 944
rect 142896 892 142948 944
rect 106188 824 106240 876
rect 123668 824 123720 876
rect 123852 824 123904 876
rect 153108 824 153160 876
rect 87144 756 87196 808
rect 110420 756 110472 808
rect 128360 756 128412 808
rect 144920 756 144972 808
rect 84844 688 84896 740
rect 276020 688 276072 740
rect 78772 552 78824 604
rect 237380 552 237432 604
rect 100760 484 100812 536
rect 218244 484 218296 536
rect 117872 416 117924 468
rect 136272 416 136324 468
rect 149060 212 149112 264
rect 256700 212 256752 264
rect 158720 144 158772 196
rect 295708 144 295760 196
rect 79324 76 79376 128
rect 253664 76 253716 128
rect 67548 8 67600 60
rect 126612 8 126664 60
rect 130292 8 130344 60
rect 143356 8 143408 60
rect 178040 8 178092 60
rect 356520 8 356572 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700670 8156 703520
rect 24320 700738 24348 703520
rect 24308 700732 24360 700738
rect 24308 700674 24360 700680
rect 8116 700664 8168 700670
rect 8116 700606 8168 700612
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 40052 496126 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 699718 73016 703520
rect 89180 700874 89208 703520
rect 89168 700868 89220 700874
rect 89168 700810 89220 700816
rect 96620 700868 96672 700874
rect 96620 700810 96672 700816
rect 95884 700800 95936 700806
rect 95884 700742 95936 700748
rect 87052 700596 87104 700602
rect 87052 700538 87104 700544
rect 84200 700528 84252 700534
rect 84200 700470 84252 700476
rect 80060 700460 80112 700466
rect 80060 700402 80112 700408
rect 77300 700392 77352 700398
rect 77300 700334 77352 700340
rect 74540 700324 74592 700330
rect 74540 700266 74592 700272
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 72424 696992 72476 696998
rect 72424 696934 72476 696940
rect 70492 683188 70544 683194
rect 70492 683130 70544 683136
rect 66260 643136 66312 643142
rect 66260 643078 66312 643084
rect 64972 616888 65024 616894
rect 64972 616830 65024 616836
rect 63500 590708 63552 590714
rect 63500 590650 63552 590656
rect 62120 563100 62172 563106
rect 62120 563042 62172 563048
rect 59452 536852 59504 536858
rect 59452 536794 59504 536800
rect 57980 510672 58032 510678
rect 57980 510614 58032 510620
rect 40040 496120 40092 496126
rect 40040 496062 40092 496068
rect 56600 484424 56652 484430
rect 56600 484366 56652 484372
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 55220 456816 55272 456822
rect 55220 456758 55272 456764
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 52460 430636 52512 430642
rect 52460 430578 52512 430584
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 35164 422340 35216 422346
rect 35164 422282 35216 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 240174 3464 241023
rect 3424 240168 3476 240174
rect 3424 240110 3476 240116
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3436 201550 3464 201855
rect 3424 201544 3476 201550
rect 3424 201486 3476 201492
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3436 187746 3464 188799
rect 3424 187740 3476 187746
rect 3424 187682 3476 187688
rect 3424 162920 3476 162926
rect 3422 162888 3424 162897
rect 3476 162888 3478 162897
rect 3422 162823 3478 162832
rect 33784 162376 33836 162382
rect 33784 162318 33836 162324
rect 20628 162308 20680 162314
rect 20628 162250 20680 162256
rect 2872 162240 2924 162246
rect 2872 162182 2924 162188
rect 1216 162172 1268 162178
rect 1216 162114 1268 162120
rect 940 159180 992 159186
rect 940 159122 992 159128
rect 848 153196 900 153202
rect 848 153138 900 153144
rect 860 17406 888 153138
rect 848 17400 900 17406
rect 848 17342 900 17348
rect 952 16658 980 159122
rect 1032 158840 1084 158846
rect 1032 158782 1084 158788
rect 940 16652 992 16658
rect 940 16594 992 16600
rect 1044 14550 1072 158782
rect 1124 157956 1176 157962
rect 1124 157898 1176 157904
rect 1032 14544 1084 14550
rect 1032 14486 1084 14492
rect 1136 11762 1164 157898
rect 1228 12374 1256 162114
rect 2780 161696 2832 161702
rect 2780 161638 2832 161644
rect 2688 160812 2740 160818
rect 2688 160754 2740 160760
rect 2412 160472 2464 160478
rect 2412 160414 2464 160420
rect 2320 158908 2372 158914
rect 2320 158850 2372 158856
rect 1308 158772 1360 158778
rect 1308 158714 1360 158720
rect 1216 12368 1268 12374
rect 1216 12310 1268 12316
rect 1124 11756 1176 11762
rect 1124 11698 1176 11704
rect 1320 6322 1348 158714
rect 2228 153332 2280 153338
rect 2228 153274 2280 153280
rect 2240 17474 2268 153274
rect 2228 17468 2280 17474
rect 2228 17410 2280 17416
rect 2332 17202 2360 158850
rect 2424 18630 2452 160414
rect 2596 160132 2648 160138
rect 2596 160074 2648 160080
rect 2504 156052 2556 156058
rect 2504 155994 2556 156000
rect 2412 18624 2464 18630
rect 2412 18566 2464 18572
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2516 14958 2544 155994
rect 2608 15026 2636 160074
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2700 12306 2728 160754
rect 2792 158778 2820 161638
rect 2884 158846 2912 162182
rect 3332 162104 3384 162110
rect 3332 162046 3384 162052
rect 2872 158840 2924 158846
rect 2872 158782 2924 158788
rect 2780 158772 2832 158778
rect 2780 158714 2832 158720
rect 3240 153740 3292 153746
rect 3240 153682 3292 153688
rect 3252 142154 3280 153682
rect 3344 153202 3372 162046
rect 17040 162036 17092 162042
rect 17040 161978 17092 161984
rect 12716 161968 12768 161974
rect 12716 161910 12768 161916
rect 4068 161900 4120 161906
rect 4068 161842 4120 161848
rect 3976 160676 4028 160682
rect 3976 160618 4028 160624
rect 3700 160608 3752 160614
rect 3700 160550 3752 160556
rect 3608 156664 3660 156670
rect 3608 156606 3660 156612
rect 3332 153196 3384 153202
rect 3332 153138 3384 153144
rect 3424 152176 3476 152182
rect 3424 152118 3476 152124
rect 3436 151814 3464 152118
rect 3436 151786 3556 151814
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3252 142126 3464 142154
rect 3436 110673 3464 142126
rect 3528 136785 3556 151786
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 135856 3568 135862
rect 3516 135798 3568 135804
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3148 97980 3200 97986
rect 3148 97922 3200 97928
rect 3160 97617 3188 97922
rect 3146 97608 3202 97617
rect 3146 97543 3202 97552
rect 2964 85536 3016 85542
rect 2964 85478 3016 85484
rect 2976 84697 3004 85478
rect 2962 84688 3018 84697
rect 2962 84623 3018 84632
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 3476 71632 3478 71641
rect 3422 71567 3478 71576
rect 3332 59356 3384 59362
rect 3332 59298 3384 59304
rect 3344 58585 3372 59298
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 32632 3476 32638
rect 3424 32574 3476 32580
rect 3436 32473 3464 32574
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3160 19417 3188 19994
rect 3146 19408 3202 19417
rect 3146 19343 3202 19352
rect 3528 17746 3556 135798
rect 3620 19922 3648 156606
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 480 1716 2926
rect 2884 480 2912 14418
rect 3436 2990 3464 15846
rect 3712 14890 3740 160550
rect 3792 160268 3844 160274
rect 3792 160210 3844 160216
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3804 14822 3832 160210
rect 3884 160200 3936 160206
rect 3884 160142 3936 160148
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3896 13122 3924 160142
rect 3988 13734 4016 160618
rect 4080 15162 4108 161842
rect 8300 161832 8352 161838
rect 8300 161774 8352 161780
rect 7656 161560 7708 161566
rect 7656 161502 7708 161508
rect 5080 159724 5132 159730
rect 5080 159666 5132 159672
rect 4804 155848 4856 155854
rect 4804 155790 4856 155796
rect 4816 20058 4844 155790
rect 4988 152584 5040 152590
rect 4988 152526 5040 152532
rect 4896 152516 4948 152522
rect 4896 152458 4948 152464
rect 4908 135862 4936 152458
rect 4896 135856 4948 135862
rect 4896 135798 4948 135804
rect 4896 134632 4948 134638
rect 4896 134574 4948 134580
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3884 13116 3936 13122
rect 3884 13058 3936 13064
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3528 6497 3556 6802
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 4172 3482 4200 7686
rect 4816 3534 4844 15982
rect 4908 14686 4936 134574
rect 5000 18698 5028 152526
rect 5092 18766 5120 159666
rect 6828 159588 6880 159594
rect 6828 159530 6880 159536
rect 6736 159384 6788 159390
rect 6736 159326 6788 159332
rect 6644 159316 6696 159322
rect 6644 159258 6696 159264
rect 6552 159248 6604 159254
rect 6552 159190 6604 159196
rect 5448 158840 5500 158846
rect 5448 158782 5500 158788
rect 5356 158772 5408 158778
rect 5356 158714 5408 158720
rect 5172 158024 5224 158030
rect 5172 157966 5224 157972
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 5184 15978 5212 157966
rect 5264 156800 5316 156806
rect 5264 156742 5316 156748
rect 5172 15972 5224 15978
rect 5172 15914 5224 15920
rect 4896 14680 4948 14686
rect 4896 14622 4948 14628
rect 5276 14618 5304 156742
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5368 13802 5396 158714
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5460 10606 5488 158782
rect 6184 158160 6236 158166
rect 6184 158102 6236 158108
rect 6196 134638 6224 158102
rect 6460 153264 6512 153270
rect 6460 153206 6512 153212
rect 6368 149116 6420 149122
rect 6368 149058 6420 149064
rect 6184 134632 6236 134638
rect 6184 134574 6236 134580
rect 6380 19990 6408 149058
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 4080 3454 4200 3482
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5264 3460 5316 3466
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 4080 480 4108 3454
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16934
rect 6472 16318 6500 153206
rect 6564 18902 6592 159190
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6656 17814 6684 159258
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6748 16386 6776 159326
rect 6736 16380 6788 16386
rect 6736 16322 6788 16328
rect 6460 16312 6512 16318
rect 6460 16254 6512 16260
rect 6840 12170 6868 159530
rect 7564 153808 7616 153814
rect 7564 153750 7616 153756
rect 7576 71670 7604 153750
rect 7668 153338 7696 161502
rect 8312 158914 8340 161774
rect 8392 161764 8444 161770
rect 8392 161706 8444 161712
rect 8300 158908 8352 158914
rect 8300 158850 8352 158856
rect 8404 157962 8432 161706
rect 12348 160948 12400 160954
rect 12348 160890 12400 160896
rect 9126 160168 9182 160177
rect 9126 160103 9182 160112
rect 8392 157956 8444 157962
rect 8392 157898 8444 157904
rect 7840 157684 7892 157690
rect 7840 157626 7892 157632
rect 7748 155372 7800 155378
rect 7748 155314 7800 155320
rect 7656 153332 7708 153338
rect 7656 153274 7708 153280
rect 7656 150476 7708 150482
rect 7656 150418 7708 150424
rect 7564 71664 7616 71670
rect 7564 71606 7616 71612
rect 7668 17542 7696 150418
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7760 17066 7788 155314
rect 7852 18222 7880 157626
rect 7932 156732 7984 156738
rect 7932 156674 7984 156680
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7944 16590 7972 156674
rect 8116 154624 8168 154630
rect 8116 154566 8168 154572
rect 8024 152652 8076 152658
rect 8024 152594 8076 152600
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 7668 480 7696 16050
rect 8036 12442 8064 152594
rect 8128 15094 8156 154566
rect 8300 154556 8352 154562
rect 8300 154498 8352 154504
rect 8208 153876 8260 153882
rect 8208 153818 8260 153824
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8220 12646 8248 153818
rect 8312 149122 8340 154498
rect 8944 154284 8996 154290
rect 8944 154226 8996 154232
rect 8300 149116 8352 149122
rect 8300 149058 8352 149064
rect 8956 32638 8984 154226
rect 9036 150544 9088 150550
rect 9036 150486 9088 150492
rect 8944 32632 8996 32638
rect 8944 32574 8996 32580
rect 9048 17202 9076 150486
rect 9140 150482 9168 160103
rect 9404 159520 9456 159526
rect 9404 159462 9456 159468
rect 9312 157956 9364 157962
rect 9312 157898 9364 157904
rect 9220 154148 9272 154154
rect 9220 154090 9272 154096
rect 9128 150476 9180 150482
rect 9128 150418 9180 150424
rect 9128 149116 9180 149122
rect 9128 149058 9180 149064
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8404 11966 8432 16594
rect 8392 11960 8444 11966
rect 8392 11902 8444 11908
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8772 480 8800 11834
rect 8956 8294 8984 17138
rect 9140 14414 9168 149058
rect 9232 17610 9260 154090
rect 9324 151814 9352 157898
rect 9416 153270 9444 159462
rect 11980 159452 12032 159458
rect 11980 159394 12032 159400
rect 9680 158092 9732 158098
rect 9680 158034 9732 158040
rect 9496 157412 9548 157418
rect 9496 157354 9548 157360
rect 9404 153264 9456 153270
rect 9404 153206 9456 153212
rect 9324 151786 9444 151814
rect 9312 150476 9364 150482
rect 9312 150418 9364 150424
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9324 12986 9352 150418
rect 9416 17882 9444 151786
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9508 15201 9536 157354
rect 9588 154692 9640 154698
rect 9588 154634 9640 154640
rect 9494 15192 9550 15201
rect 9494 15127 9550 15136
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9600 10334 9628 154634
rect 9692 154630 9720 158034
rect 10048 157616 10100 157622
rect 10048 157558 10100 157564
rect 9680 154624 9732 154630
rect 9680 154566 9732 154572
rect 10060 154154 10088 157558
rect 10968 156596 11020 156602
rect 10968 156538 11020 156544
rect 10784 156392 10836 156398
rect 10784 156334 10836 156340
rect 10232 155984 10284 155990
rect 10232 155926 10284 155932
rect 10048 154148 10100 154154
rect 10048 154090 10100 154096
rect 10244 149122 10272 155926
rect 10324 155916 10376 155922
rect 10324 155858 10376 155864
rect 10232 149116 10284 149122
rect 10232 149058 10284 149064
rect 10336 59362 10364 155858
rect 10416 154216 10468 154222
rect 10416 154158 10468 154164
rect 10324 59356 10376 59362
rect 10324 59298 10376 59304
rect 10324 56976 10376 56982
rect 10324 56918 10376 56924
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9588 10328 9640 10334
rect 9588 10270 9640 10276
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 17274
rect 10336 13530 10364 56918
rect 10428 19786 10456 154158
rect 10692 151904 10744 151910
rect 10506 151872 10562 151881
rect 10692 151846 10744 151852
rect 10506 151807 10562 151816
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10520 18358 10548 151807
rect 10600 150612 10652 150618
rect 10600 150554 10652 150560
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10612 17950 10640 150554
rect 10600 17944 10652 17950
rect 10600 17886 10652 17892
rect 10704 17762 10732 151846
rect 10612 17734 10732 17762
rect 10612 16454 10640 17734
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10612 12102 10640 14962
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10704 12034 10732 17478
rect 10796 17134 10824 156334
rect 10876 154624 10928 154630
rect 10876 154566 10928 154572
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10888 16522 10916 154566
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10692 12028 10744 12034
rect 10692 11970 10744 11976
rect 10796 9926 10824 15098
rect 10980 15026 11008 156538
rect 11888 155576 11940 155582
rect 11888 155518 11940 155524
rect 11796 152040 11848 152046
rect 11796 151982 11848 151988
rect 11704 151972 11756 151978
rect 11704 151914 11756 151920
rect 11716 56982 11744 151914
rect 11704 56976 11756 56982
rect 11704 56918 11756 56924
rect 11808 18834 11836 151982
rect 11900 20058 11928 155518
rect 11992 150550 12020 159394
rect 12256 155440 12308 155446
rect 12256 155382 12308 155388
rect 12072 155100 12124 155106
rect 12072 155042 12124 155048
rect 11980 150544 12032 150550
rect 11980 150486 12032 150492
rect 11980 147688 12032 147694
rect 11980 147630 12032 147636
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10888 11082 10916 14894
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10980 9625 11008 13738
rect 11072 10470 11100 16526
rect 11992 13054 12020 147630
rect 12084 19174 12112 155042
rect 12164 154148 12216 154154
rect 12164 154090 12216 154096
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12176 17814 12204 154090
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12268 17746 12296 155382
rect 12360 154562 12388 160890
rect 12532 160880 12584 160886
rect 12532 160822 12584 160828
rect 12440 156120 12492 156126
rect 12440 156062 12492 156068
rect 12348 154556 12400 154562
rect 12348 154498 12400 154504
rect 12452 151814 12480 156062
rect 12544 152522 12572 160822
rect 12728 159594 12756 161910
rect 15844 161628 15896 161634
rect 15844 161570 15896 161576
rect 13268 160336 13320 160342
rect 13268 160278 13320 160284
rect 12716 159588 12768 159594
rect 12716 159530 12768 159536
rect 12624 158908 12676 158914
rect 12624 158850 12676 158856
rect 12636 155378 12664 158850
rect 12992 157480 13044 157486
rect 12992 157422 13044 157428
rect 12900 156256 12952 156262
rect 12900 156198 12952 156204
rect 12624 155372 12676 155378
rect 12624 155314 12676 155320
rect 12532 152516 12584 152522
rect 12532 152458 12584 152464
rect 12360 151786 12480 151814
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11980 13048 12032 13054
rect 12360 13025 12388 151786
rect 12912 150482 12940 156198
rect 13004 154698 13032 157422
rect 13280 155990 13308 160278
rect 14280 158976 14332 158982
rect 14280 158918 14332 158924
rect 13728 157888 13780 157894
rect 13728 157830 13780 157836
rect 13268 155984 13320 155990
rect 13268 155926 13320 155932
rect 13360 155984 13412 155990
rect 13360 155926 13412 155932
rect 13268 155644 13320 155650
rect 13268 155586 13320 155592
rect 12992 154692 13044 154698
rect 12992 154634 13044 154640
rect 12992 152244 13044 152250
rect 12992 152186 13044 152192
rect 12900 150476 12952 150482
rect 12900 150418 12952 150424
rect 13004 85542 13032 152186
rect 13176 151768 13228 151774
rect 13176 151710 13228 151716
rect 13084 150476 13136 150482
rect 13084 150418 13136 150424
rect 12992 85536 13044 85542
rect 12992 85478 13044 85484
rect 12992 82884 13044 82890
rect 12992 82826 13044 82832
rect 13004 20534 13032 82826
rect 13096 20602 13124 150418
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 13188 16697 13216 151710
rect 13280 20126 13308 155586
rect 13268 20120 13320 20126
rect 13268 20062 13320 20068
rect 13372 18630 13400 155926
rect 13452 155508 13504 155514
rect 13452 155450 13504 155456
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13268 17944 13320 17950
rect 13268 17886 13320 17892
rect 13174 16688 13230 16697
rect 13174 16623 13230 16632
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 11980 12990 12032 12996
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 12452 9654 12480 12106
rect 12440 9648 12492 9654
rect 10966 9616 11022 9625
rect 12440 9590 12492 9596
rect 10966 9551 11022 9560
rect 11152 4888 11204 4894
rect 11152 4830 11204 4836
rect 11164 480 11192 4830
rect 13096 3534 13124 16118
rect 13280 10402 13308 17886
rect 13464 17882 13492 155450
rect 13634 153776 13690 153785
rect 13634 153711 13690 153720
rect 13542 153232 13598 153241
rect 13542 153167 13598 153176
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13372 15162 13400 17818
rect 13452 17400 13504 17406
rect 13452 17342 13504 17348
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13464 11150 13492 17342
rect 13556 15774 13584 153167
rect 13544 15768 13596 15774
rect 13544 15710 13596 15716
rect 13648 13258 13676 153711
rect 13740 15842 13768 157830
rect 14292 147694 14320 158918
rect 15016 157548 15068 157554
rect 15016 157490 15068 157496
rect 14462 156088 14518 156097
rect 14462 156023 14518 156032
rect 14372 155032 14424 155038
rect 14372 154974 14424 154980
rect 14280 147688 14332 147694
rect 14280 147630 14332 147636
rect 14384 45558 14412 154974
rect 14476 150482 14504 156023
rect 14648 154760 14700 154766
rect 14648 154702 14700 154708
rect 14830 154728 14886 154737
rect 14554 153368 14610 153377
rect 14554 153303 14610 153312
rect 14464 150476 14516 150482
rect 14464 150418 14516 150424
rect 14464 149116 14516 149122
rect 14464 149058 14516 149064
rect 14372 45552 14424 45558
rect 14372 45494 14424 45500
rect 14476 18018 14504 149058
rect 14568 18086 14596 153303
rect 14660 18154 14688 154702
rect 14830 154663 14886 154672
rect 14738 154184 14794 154193
rect 14738 154119 14794 154128
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14464 18012 14516 18018
rect 14464 17954 14516 17960
rect 14752 15881 14780 154119
rect 14844 16561 14872 154663
rect 14924 152788 14976 152794
rect 14924 152730 14976 152736
rect 14830 16552 14886 16561
rect 14830 16487 14886 16496
rect 14738 15872 14794 15881
rect 13728 15836 13780 15842
rect 14738 15807 14794 15816
rect 13728 15778 13780 15784
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13832 13734 13860 14486
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 14936 10674 14964 152730
rect 15028 14521 15056 157490
rect 15856 153202 15884 161570
rect 16672 159588 16724 159594
rect 16672 159530 16724 159536
rect 16488 156528 16540 156534
rect 16488 156470 16540 156476
rect 16396 155780 16448 155786
rect 16396 155722 16448 155728
rect 15936 155712 15988 155718
rect 15936 155654 15988 155660
rect 15108 153196 15160 153202
rect 15108 153138 15160 153144
rect 15844 153196 15896 153202
rect 15844 153138 15896 153144
rect 15014 14512 15070 14521
rect 15014 14447 15070 14456
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 13268 10396 13320 10402
rect 13268 10338 13320 10344
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12360 480 12388 3470
rect 13556 480 13584 9114
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 10474
rect 15120 7682 15148 153138
rect 15752 152516 15804 152522
rect 15752 152458 15804 152464
rect 15764 149122 15792 152458
rect 15948 150618 15976 155654
rect 16304 154692 16356 154698
rect 16304 154634 16356 154640
rect 16028 152992 16080 152998
rect 16028 152934 16080 152940
rect 15936 150612 15988 150618
rect 15936 150554 15988 150560
rect 15936 149728 15988 149734
rect 15936 149670 15988 149676
rect 15752 149116 15804 149122
rect 15752 149058 15804 149064
rect 15948 20670 15976 149670
rect 15936 20664 15988 20670
rect 15936 20606 15988 20612
rect 16040 19961 16068 152934
rect 16212 152924 16264 152930
rect 16212 152866 16264 152872
rect 16120 151088 16172 151094
rect 16120 151030 16172 151036
rect 16026 19952 16082 19961
rect 16026 19887 16082 19896
rect 15660 18896 15712 18902
rect 15660 18838 15712 18844
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15212 16250 15240 18634
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15396 15638 15424 18702
rect 15568 17400 15620 17406
rect 15568 17342 15620 17348
rect 15476 16380 15528 16386
rect 15476 16322 15528 16328
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15396 14890 15424 15030
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15212 8974 15240 11698
rect 15304 11490 15332 14826
rect 15488 13666 15516 16322
rect 15476 13660 15528 13666
rect 15476 13602 15528 13608
rect 15292 11484 15344 11490
rect 15292 11426 15344 11432
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15108 7676 15160 7682
rect 15108 7618 15160 7624
rect 15580 6914 15608 17342
rect 15672 14346 15700 18838
rect 16132 18698 16160 151030
rect 16224 18902 16252 152866
rect 16316 19650 16344 154634
rect 16304 19644 16356 19650
rect 16304 19586 16356 19592
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16408 18290 16436 155722
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16500 16522 16528 156470
rect 16684 152590 16712 159530
rect 16672 152584 16724 152590
rect 16672 152526 16724 152532
rect 17052 149734 17080 161978
rect 20260 160404 20312 160410
rect 20260 160346 20312 160352
rect 18420 159656 18472 159662
rect 18420 159598 18472 159604
rect 18050 159352 18106 159361
rect 18050 159287 18106 159296
rect 17408 157820 17460 157826
rect 17408 157762 17460 157768
rect 17224 154964 17276 154970
rect 17224 154906 17276 154912
rect 17132 153196 17184 153202
rect 17132 153138 17184 153144
rect 17040 149728 17092 149734
rect 17040 149670 17092 149676
rect 17144 82890 17172 153138
rect 17132 82884 17184 82890
rect 17132 82826 17184 82832
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 17052 19718 17080 27066
rect 17236 22094 17264 154906
rect 17420 152658 17448 157762
rect 17868 157752 17920 157758
rect 17868 157694 17920 157700
rect 17776 156460 17828 156466
rect 17776 156402 17828 156408
rect 17684 153672 17736 153678
rect 17684 153614 17736 153620
rect 17500 153604 17552 153610
rect 17500 153546 17552 153552
rect 17408 152652 17460 152658
rect 17408 152594 17460 152600
rect 17316 150544 17368 150550
rect 17316 150486 17368 150492
rect 17328 27130 17356 150486
rect 17408 150476 17460 150482
rect 17408 150418 17460 150424
rect 17316 27124 17368 27130
rect 17316 27066 17368 27072
rect 17420 27010 17448 150418
rect 17144 22066 17264 22094
rect 17328 26982 17448 27010
rect 17144 21434 17172 22066
rect 17144 21406 17264 21434
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16764 18012 16816 18018
rect 16764 17954 16816 17960
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 15752 15836 15804 15842
rect 15752 15778 15804 15784
rect 15764 14958 15792 15778
rect 16776 15230 16804 17954
rect 16764 15224 16816 15230
rect 16764 15166 16816 15172
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 16960 13190 16988 18022
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 15580 6886 15976 6914
rect 15948 480 15976 6886
rect 17052 480 17080 14486
rect 17144 9314 17172 20470
rect 17132 9308 17184 9314
rect 17132 9250 17184 9256
rect 17236 6866 17264 21406
rect 17328 18562 17356 26982
rect 17512 26874 17540 153546
rect 17592 153536 17644 153542
rect 17592 153478 17644 153484
rect 17420 26846 17540 26874
rect 17420 18601 17448 26846
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17512 18766 17540 26726
rect 17604 19310 17632 153478
rect 17696 26790 17724 153614
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17500 18760 17552 18766
rect 17696 18737 17724 20538
rect 17788 19854 17816 156402
rect 17880 153882 17908 157694
rect 18064 155650 18092 159287
rect 18234 157448 18290 157457
rect 18234 157383 18290 157392
rect 18052 155644 18104 155650
rect 18052 155586 18104 155592
rect 17868 153876 17920 153882
rect 17868 153818 17920 153824
rect 18144 153876 18196 153882
rect 18144 153818 18196 153824
rect 17868 153264 17920 153270
rect 17868 153206 17920 153212
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17500 18702 17552 18708
rect 17682 18728 17738 18737
rect 17682 18663 17738 18672
rect 17684 18624 17736 18630
rect 17406 18592 17462 18601
rect 17316 18556 17368 18562
rect 17684 18566 17736 18572
rect 17406 18527 17462 18536
rect 17316 18498 17368 18504
rect 17696 17785 17724 18566
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17682 17776 17738 17785
rect 17682 17711 17738 17720
rect 17788 16930 17816 18090
rect 17776 16924 17828 16930
rect 17776 16866 17828 16872
rect 17880 15842 17908 153206
rect 18156 152046 18184 153818
rect 18144 152040 18196 152046
rect 18144 151982 18196 151988
rect 18248 151842 18276 157383
rect 18328 155304 18380 155310
rect 18328 155246 18380 155252
rect 18236 151836 18288 151842
rect 18236 151778 18288 151784
rect 18340 150414 18368 155246
rect 18432 151978 18460 159598
rect 18788 159044 18840 159050
rect 18788 158986 18840 158992
rect 18800 155718 18828 158986
rect 19248 156868 19300 156874
rect 19248 156810 19300 156816
rect 19064 156188 19116 156194
rect 19064 156130 19116 156136
rect 18788 155712 18840 155718
rect 18788 155654 18840 155660
rect 18512 155168 18564 155174
rect 18512 155110 18564 155116
rect 18420 151972 18472 151978
rect 18420 151914 18472 151920
rect 18328 150408 18380 150414
rect 18328 150350 18380 150356
rect 18524 97986 18552 155110
rect 18788 153400 18840 153406
rect 18788 153342 18840 153348
rect 18696 153332 18748 153338
rect 18696 153274 18748 153280
rect 18604 152108 18656 152114
rect 18604 152050 18656 152056
rect 18512 97980 18564 97986
rect 18512 97922 18564 97928
rect 18512 20664 18564 20670
rect 18512 20606 18564 20612
rect 18052 18488 18104 18494
rect 18052 18430 18104 18436
rect 17868 15836 17920 15842
rect 17868 15778 17920 15784
rect 18064 15298 18092 18430
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18144 17468 18196 17474
rect 18144 17410 18196 17416
rect 18052 15292 18104 15298
rect 18052 15234 18104 15240
rect 18156 13870 18184 17410
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18248 13598 18276 17614
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18236 13592 18288 13598
rect 18236 13534 18288 13540
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17696 3466 17724 6326
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 13262
rect 18432 11694 18460 17002
rect 18524 15570 18552 20606
rect 18616 19242 18644 152050
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18708 18630 18736 153274
rect 18800 19038 18828 153342
rect 18880 152312 18932 152318
rect 18880 152254 18932 152260
rect 18788 19032 18840 19038
rect 18788 18974 18840 18980
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18892 17921 18920 152254
rect 18972 152040 19024 152046
rect 18972 151982 19024 151988
rect 18878 17912 18934 17921
rect 18878 17847 18934 17856
rect 18984 17241 19012 151982
rect 19076 20670 19104 156130
rect 19154 155000 19210 155009
rect 19154 154935 19210 154944
rect 19064 20664 19116 20670
rect 19064 20606 19116 20612
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18970 17232 19026 17241
rect 18970 17167 19026 17176
rect 18694 16688 18750 16697
rect 18694 16623 18750 16632
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18604 14680 18656 14686
rect 18604 14622 18656 14628
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18616 9450 18644 14622
rect 18708 11762 18736 16623
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18788 11960 18840 11966
rect 18788 11902 18840 11908
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18800 9518 18828 11902
rect 18892 11558 18920 14894
rect 18984 13938 19012 16458
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 19076 11966 19104 18838
rect 19168 18494 19196 154935
rect 19156 18488 19208 18494
rect 19156 18430 19208 18436
rect 19260 16574 19288 156810
rect 20168 156324 20220 156330
rect 20168 156266 20220 156272
rect 19706 155136 19762 155145
rect 19706 155071 19762 155080
rect 19616 154556 19668 154562
rect 19616 154498 19668 154504
rect 19628 150550 19656 154498
rect 19616 150544 19668 150550
rect 19616 150486 19668 150492
rect 19720 150482 19748 155071
rect 19798 154864 19854 154873
rect 19798 154799 19854 154808
rect 19812 151094 19840 154799
rect 19892 153128 19944 153134
rect 19892 153070 19944 153076
rect 19904 151910 19932 153070
rect 19984 151972 20036 151978
rect 19984 151914 20036 151920
rect 19892 151904 19944 151910
rect 19892 151846 19944 151852
rect 19800 151088 19852 151094
rect 19800 151030 19852 151036
rect 19708 150476 19760 150482
rect 19708 150418 19760 150424
rect 19800 20664 19852 20670
rect 19800 20606 19852 20612
rect 19708 20120 19760 20126
rect 19708 20062 19760 20068
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19340 17468 19392 17474
rect 19340 17410 19392 17416
rect 19168 16546 19288 16574
rect 19352 16574 19380 17410
rect 19352 16546 19472 16574
rect 19168 14958 19196 16546
rect 19248 16312 19300 16318
rect 19248 16254 19300 16260
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 12345 19196 14758
rect 19260 14754 19288 16254
rect 19248 14748 19300 14754
rect 19248 14690 19300 14696
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19154 12336 19210 12345
rect 19154 12271 19210 12280
rect 19064 11960 19116 11966
rect 19064 11902 19116 11908
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 19352 10742 19380 13806
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 19444 480 19472 16546
rect 19628 15502 19656 19994
rect 19720 19281 19748 20062
rect 19706 19272 19762 19281
rect 19706 19207 19762 19216
rect 19812 18970 19840 20606
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19904 14686 19932 19926
rect 19996 17950 20024 151914
rect 20076 151904 20128 151910
rect 20076 151846 20128 151852
rect 19984 17944 20036 17950
rect 19984 17886 20036 17892
rect 20088 16862 20116 151846
rect 20076 16856 20128 16862
rect 20076 16798 20128 16804
rect 20180 16289 20208 156266
rect 20166 16280 20222 16289
rect 20166 16215 20222 16224
rect 20168 15292 20220 15298
rect 20168 15234 20220 15240
rect 19892 14680 19944 14686
rect 19892 14622 19944 14628
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19628 9110 19656 12038
rect 20180 11626 20208 15234
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20272 9246 20300 160346
rect 20640 159730 20668 162250
rect 20628 159724 20680 159730
rect 20628 159666 20680 159672
rect 33796 159662 33824 162318
rect 35176 160750 35204 422282
rect 49700 378208 49752 378214
rect 49700 378150 49752 378156
rect 48412 351960 48464 351966
rect 48412 351902 48464 351908
rect 46940 324352 46992 324358
rect 46940 324294 46992 324300
rect 45560 298172 45612 298178
rect 45560 298114 45612 298120
rect 42892 271924 42944 271930
rect 42892 271866 42944 271872
rect 41420 244316 41472 244322
rect 41420 244258 41472 244264
rect 40040 231872 40092 231878
rect 40040 231814 40092 231820
rect 38660 205692 38712 205698
rect 38660 205634 38712 205640
rect 35900 191888 35952 191894
rect 35900 191830 35952 191836
rect 35164 160744 35216 160750
rect 35164 160686 35216 160692
rect 33784 159656 33836 159662
rect 33784 159598 33836 159604
rect 20626 158808 20682 158817
rect 20626 158743 20682 158752
rect 20352 158228 20404 158234
rect 20352 158170 20404 158176
rect 20364 153202 20392 158170
rect 20352 153196 20404 153202
rect 20352 153138 20404 153144
rect 20640 152998 20668 158743
rect 21364 155712 21416 155718
rect 21364 155654 21416 155660
rect 20904 155644 20956 155650
rect 20904 155586 20956 155592
rect 20628 152992 20680 152998
rect 20628 152934 20680 152940
rect 20916 152794 20944 155586
rect 21376 152930 21404 155654
rect 23480 155576 23532 155582
rect 23480 155518 23532 155524
rect 22098 155408 22154 155417
rect 22098 155343 22154 155352
rect 22112 153785 22140 155343
rect 22192 154692 22244 154698
rect 22192 154634 22244 154640
rect 22098 153776 22154 153785
rect 22098 153711 22154 153720
rect 22204 153649 22232 154634
rect 23492 153950 23520 155518
rect 28816 155508 28868 155514
rect 28816 155450 28868 155456
rect 26240 154828 26292 154834
rect 26240 154770 26292 154776
rect 26252 154630 26280 154770
rect 27528 154760 27580 154766
rect 27528 154702 27580 154708
rect 26240 154624 26292 154630
rect 26240 154566 26292 154572
rect 23480 153944 23532 153950
rect 23480 153886 23532 153892
rect 26146 153776 26202 153785
rect 26146 153711 26202 153720
rect 22190 153640 22246 153649
rect 22190 153575 22246 153584
rect 24306 153504 24362 153513
rect 23204 153468 23256 153474
rect 24306 153439 24362 153448
rect 23204 153410 23256 153416
rect 21364 152924 21416 152930
rect 21364 152866 21416 152872
rect 20904 152788 20956 152794
rect 20904 152730 20956 152736
rect 23216 152674 23244 153410
rect 24320 152674 24348 153439
rect 25410 152688 25466 152697
rect 22908 152646 23244 152674
rect 24012 152646 24348 152674
rect 25116 152646 25410 152674
rect 26160 152674 26188 153711
rect 27540 153202 27568 154702
rect 28722 154592 28778 154601
rect 28722 154527 28778 154536
rect 27528 153196 27580 153202
rect 27528 153138 27580 153144
rect 28736 152674 28764 154527
rect 28828 153134 28856 155450
rect 35622 155408 35678 155417
rect 35256 155372 35308 155378
rect 35622 155343 35678 155352
rect 35256 155314 35308 155320
rect 31666 155272 31722 155281
rect 31666 155207 31722 155216
rect 34152 155236 34204 155242
rect 31024 154828 31076 154834
rect 31024 154770 31076 154776
rect 30196 154692 30248 154698
rect 30196 154634 30248 154640
rect 28908 154624 28960 154630
rect 28908 154566 28960 154572
rect 28920 154465 28948 154566
rect 28906 154456 28962 154465
rect 28906 154391 28962 154400
rect 29826 153912 29882 153921
rect 29826 153847 29882 153856
rect 28816 153128 28868 153134
rect 28816 153070 28868 153076
rect 29840 152674 29868 153847
rect 30208 153066 30236 154634
rect 30288 154148 30340 154154
rect 30288 154090 30340 154096
rect 30196 153060 30248 153066
rect 30196 153002 30248 153008
rect 30300 152998 30328 154090
rect 30932 154080 30984 154086
rect 30932 154022 30984 154028
rect 30838 153640 30894 153649
rect 30838 153575 30894 153584
rect 30288 152992 30340 152998
rect 30288 152934 30340 152940
rect 30852 152674 30880 153575
rect 30944 153202 30972 154022
rect 31036 153202 31064 154770
rect 30932 153196 30984 153202
rect 30932 153138 30984 153144
rect 31024 153196 31076 153202
rect 31024 153138 31076 153144
rect 26160 152646 26220 152674
rect 28428 152646 28764 152674
rect 29532 152646 29868 152674
rect 30636 152646 30880 152674
rect 31680 152674 31708 155207
rect 34152 155178 34204 155184
rect 32956 153944 33008 153950
rect 32956 153886 33008 153892
rect 33048 153944 33100 153950
rect 33048 153886 33100 153892
rect 32968 152930 32996 153886
rect 33060 153134 33088 153886
rect 34164 153882 34192 155178
rect 34428 154148 34480 154154
rect 34428 154090 34480 154096
rect 34152 153876 34204 153882
rect 34152 153818 34204 153824
rect 33048 153128 33100 153134
rect 33048 153070 33100 153076
rect 32956 152924 33008 152930
rect 32956 152866 33008 152872
rect 31680 152646 31740 152674
rect 25410 152623 25466 152632
rect 33046 152552 33102 152561
rect 32844 152510 33046 152538
rect 34440 152522 34468 154090
rect 34978 154048 35034 154057
rect 34978 153983 35034 153992
rect 34992 153474 35020 153983
rect 34980 153468 35032 153474
rect 34980 153410 35032 153416
rect 35268 152674 35296 155314
rect 35636 153882 35664 155343
rect 35912 154630 35940 191830
rect 37372 178084 37424 178090
rect 37372 178026 37424 178032
rect 37384 171134 37412 178026
rect 38672 171134 38700 205634
rect 40052 171134 40080 231814
rect 37384 171106 37964 171134
rect 38672 171106 39068 171134
rect 40052 171106 40172 171134
rect 35992 165640 36044 165646
rect 35992 165582 36044 165588
rect 35900 154624 35952 154630
rect 35900 154566 35952 154572
rect 35716 154216 35768 154222
rect 35716 154158 35768 154164
rect 35624 153876 35676 153882
rect 35624 153818 35676 153824
rect 35346 153232 35402 153241
rect 35346 153167 35402 153176
rect 35052 152646 35296 152674
rect 35360 152522 35388 153167
rect 35728 153066 35756 154158
rect 35808 154012 35860 154018
rect 35808 153954 35860 153960
rect 35820 153202 35848 153954
rect 35808 153196 35860 153202
rect 35808 153138 35860 153144
rect 35716 153060 35768 153066
rect 35716 153002 35768 153008
rect 36004 152674 36032 165582
rect 36912 154624 36964 154630
rect 36912 154566 36964 154572
rect 36924 152674 36952 154566
rect 37936 152674 37964 171106
rect 39040 152674 39068 171106
rect 40144 152674 40172 171106
rect 41432 156942 41460 244258
rect 41512 218068 41564 218074
rect 41512 218010 41564 218016
rect 41420 156936 41472 156942
rect 41420 156878 41472 156884
rect 41524 152674 41552 218010
rect 42904 171134 42932 271866
rect 44180 258120 44232 258126
rect 44180 258062 44232 258068
rect 44192 171134 44220 258062
rect 45572 171134 45600 298114
rect 42904 171106 43484 171134
rect 44192 171106 44588 171134
rect 45572 171106 45692 171134
rect 42432 156936 42484 156942
rect 42432 156878 42484 156884
rect 42444 152674 42472 156878
rect 43456 152674 43484 171106
rect 44560 152674 44588 171106
rect 45664 152674 45692 171106
rect 46952 152674 46980 324294
rect 47032 311908 47084 311914
rect 47032 311850 47084 311856
rect 47044 171134 47072 311850
rect 48424 171134 48452 351902
rect 49712 171134 49740 378150
rect 51080 364404 51132 364410
rect 51080 364346 51132 364352
rect 51092 171134 51120 364346
rect 47044 171106 47900 171134
rect 48424 171106 49004 171134
rect 49712 171106 50108 171134
rect 51092 171106 51212 171134
rect 47872 152674 47900 171106
rect 48976 152674 49004 171106
rect 50080 152674 50108 171106
rect 51184 152674 51212 171106
rect 52472 156942 52500 430578
rect 53932 418192 53984 418198
rect 53932 418134 53984 418140
rect 52552 404388 52604 404394
rect 52552 404330 52604 404336
rect 52460 156936 52512 156942
rect 52460 156878 52512 156884
rect 52564 152674 52592 404330
rect 53944 171134 53972 418134
rect 55232 171134 55260 456758
rect 56612 171134 56640 484366
rect 53944 171106 54524 171134
rect 55232 171106 55628 171134
rect 56612 171106 56732 171134
rect 53472 156936 53524 156942
rect 53472 156878 53524 156884
rect 53484 152674 53512 156878
rect 54496 152674 54524 171106
rect 55600 152674 55628 171106
rect 56704 152674 56732 171106
rect 57992 156942 58020 510614
rect 58072 470620 58124 470626
rect 58072 470562 58124 470568
rect 57980 156936 58032 156942
rect 57980 156878 58032 156884
rect 58084 152674 58112 470562
rect 59464 171134 59492 536794
rect 60740 524476 60792 524482
rect 60740 524418 60792 524424
rect 60752 171134 60780 524418
rect 62132 171134 62160 563042
rect 59464 171106 60044 171134
rect 60752 171106 61148 171134
rect 62132 171106 62252 171134
rect 58992 156936 59044 156942
rect 58992 156878 59044 156884
rect 59004 152674 59032 156878
rect 60016 152674 60044 171106
rect 61120 152674 61148 171106
rect 62224 152674 62252 171106
rect 63512 152674 63540 590650
rect 63592 576904 63644 576910
rect 63592 576846 63644 576852
rect 63604 171134 63632 576846
rect 64984 171134 65012 616830
rect 66272 171134 66300 643078
rect 67640 630692 67692 630698
rect 67640 630634 67692 630640
rect 67652 171134 67680 630634
rect 70504 171134 70532 683130
rect 63604 171106 64460 171134
rect 64984 171106 65564 171134
rect 66272 171106 66668 171134
rect 67652 171106 67772 171134
rect 70504 171106 71084 171134
rect 64432 152674 64460 171106
rect 65536 152674 65564 171106
rect 66640 152674 66668 171106
rect 67744 152674 67772 171106
rect 69664 161492 69716 161498
rect 69664 161434 69716 161440
rect 69572 161016 69624 161022
rect 69572 160958 69624 160964
rect 69584 158166 69612 160958
rect 69676 159361 69704 161434
rect 69662 159352 69718 159361
rect 69662 159287 69718 159296
rect 69664 159112 69716 159118
rect 69664 159054 69716 159060
rect 69572 158160 69624 158166
rect 69572 158102 69624 158108
rect 69570 157992 69626 158001
rect 69570 157927 69626 157936
rect 69584 152674 69612 157927
rect 69676 156806 69704 159054
rect 69664 156800 69716 156806
rect 69664 156742 69716 156748
rect 70308 156800 70360 156806
rect 70308 156742 70360 156748
rect 36004 152646 36156 152674
rect 36924 152646 37260 152674
rect 37936 152646 38364 152674
rect 39040 152646 39468 152674
rect 40144 152646 40572 152674
rect 41524 152646 41676 152674
rect 42444 152646 42780 152674
rect 43456 152646 43884 152674
rect 44560 152646 44988 152674
rect 45664 152646 46092 152674
rect 46952 152646 47196 152674
rect 47872 152646 48300 152674
rect 48976 152646 49404 152674
rect 50080 152646 50508 152674
rect 51184 152646 51612 152674
rect 52564 152646 52716 152674
rect 53484 152646 53820 152674
rect 54496 152646 54924 152674
rect 55600 152646 56028 152674
rect 56704 152646 57132 152674
rect 58084 152646 58236 152674
rect 59004 152646 59340 152674
rect 60016 152646 60444 152674
rect 61120 152646 61548 152674
rect 62224 152646 62652 152674
rect 63512 152646 63756 152674
rect 64432 152646 64860 152674
rect 65536 152646 65964 152674
rect 66640 152646 67068 152674
rect 67744 152646 68172 152674
rect 69276 152646 69612 152674
rect 70320 152674 70348 156742
rect 71056 152674 71084 171106
rect 72436 156806 72464 696934
rect 73434 162072 73490 162081
rect 73434 162007 73490 162016
rect 73252 160540 73304 160546
rect 73252 160482 73304 160488
rect 73264 158234 73292 160482
rect 73344 159656 73396 159662
rect 73344 159598 73396 159604
rect 73252 158228 73304 158234
rect 73252 158170 73304 158176
rect 73160 158160 73212 158166
rect 73160 158102 73212 158108
rect 73172 156874 73200 158102
rect 73160 156868 73212 156874
rect 73160 156810 73212 156816
rect 72424 156800 72476 156806
rect 72424 156742 72476 156748
rect 73356 156670 73384 159598
rect 73344 156664 73396 156670
rect 72882 156632 72938 156641
rect 73344 156606 73396 156612
rect 72882 156567 72938 156576
rect 72896 152674 72924 156567
rect 70320 152646 70380 152674
rect 71056 152646 71484 152674
rect 72588 152646 72924 152674
rect 73448 152674 73476 162007
rect 74552 152674 74580 700266
rect 76564 699712 76616 699718
rect 76564 699654 76616 699660
rect 76576 170406 76604 699654
rect 77312 171134 77340 700334
rect 77312 171106 77708 171134
rect 76564 170400 76616 170406
rect 76564 170342 76616 170348
rect 76564 164892 76616 164898
rect 76564 164834 76616 164840
rect 75828 156800 75880 156806
rect 75828 156742 75880 156748
rect 75840 152674 75868 156742
rect 76576 152674 76604 164834
rect 77680 152674 77708 171106
rect 78588 158228 78640 158234
rect 78588 158170 78640 158176
rect 78600 156738 78628 158170
rect 79508 156868 79560 156874
rect 79508 156810 79560 156816
rect 78588 156732 78640 156738
rect 78588 156674 78640 156680
rect 79520 152674 79548 156810
rect 80072 156738 80100 700402
rect 84212 171134 84240 700470
rect 85580 693456 85632 693462
rect 85580 693398 85632 693404
rect 85592 171134 85620 693398
rect 87064 171134 87092 700538
rect 95240 698964 95292 698970
rect 95240 698906 95292 698912
rect 92572 696244 92624 696250
rect 92572 696186 92624 696192
rect 88340 494760 88392 494766
rect 88340 494702 88392 494708
rect 88352 171134 88380 494702
rect 91100 173188 91152 173194
rect 91100 173130 91152 173136
rect 89720 171828 89772 171834
rect 89720 171770 89772 171776
rect 89732 171134 89760 171770
rect 84212 171106 84332 171134
rect 85592 171106 86540 171134
rect 87064 171106 87644 171134
rect 88352 171106 88748 171134
rect 89732 171106 89852 171134
rect 83188 169040 83240 169046
rect 83188 168982 83240 168988
rect 80152 167680 80204 167686
rect 80152 167622 80204 167628
rect 80060 156732 80112 156738
rect 80060 156674 80112 156680
rect 73448 152646 73692 152674
rect 74552 152646 74796 152674
rect 75840 152646 75900 152674
rect 76576 152646 77004 152674
rect 77680 152646 78108 152674
rect 79212 152646 79548 152674
rect 80164 152674 80192 167622
rect 82728 156800 82780 156806
rect 82728 156742 82780 156748
rect 81072 156732 81124 156738
rect 81072 156674 81124 156680
rect 81084 152674 81112 156674
rect 82740 152674 82768 156742
rect 80164 152646 80316 152674
rect 81084 152646 81420 152674
rect 82524 152646 82768 152674
rect 83200 152674 83228 168982
rect 84304 152674 84332 171106
rect 86132 156868 86184 156874
rect 86132 156810 86184 156816
rect 86144 152674 86172 156810
rect 83200 152646 83628 152674
rect 84304 152646 84732 152674
rect 85836 152646 86172 152674
rect 86512 152674 86540 171106
rect 87616 152674 87644 171106
rect 88720 152674 88748 171106
rect 89824 152674 89852 171106
rect 91112 152674 91140 173130
rect 92584 171134 92612 696186
rect 94504 397520 94556 397526
rect 94504 397462 94556 397468
rect 92584 171106 93164 171134
rect 92386 159352 92442 159361
rect 92386 159287 92442 159296
rect 92400 152674 92428 159287
rect 93136 152674 93164 171106
rect 94516 158302 94544 397462
rect 95252 171134 95280 698906
rect 95252 171106 95372 171134
rect 94504 158296 94556 158302
rect 94504 158238 94556 158244
rect 94964 155576 95016 155582
rect 94964 155518 95016 155524
rect 94320 155440 94372 155446
rect 94320 155382 94372 155388
rect 94332 154222 94360 155382
rect 94320 154216 94372 154222
rect 94320 154158 94372 154164
rect 94976 152674 95004 155518
rect 95148 154080 95200 154086
rect 95148 154022 95200 154028
rect 86512 152646 86940 152674
rect 87616 152646 88044 152674
rect 88720 152646 89148 152674
rect 89824 152646 90252 152674
rect 91112 152646 91356 152674
rect 92400 152646 92460 152674
rect 93136 152646 93564 152674
rect 94668 152646 95004 152674
rect 95160 152561 95188 154022
rect 95344 152674 95372 171106
rect 95896 155582 95924 700742
rect 96632 156942 96660 700810
rect 100760 700732 100812 700738
rect 100760 700674 100812 700680
rect 99380 700664 99432 700670
rect 99380 700606 99432 700612
rect 98092 496120 98144 496126
rect 98092 496062 98144 496068
rect 98104 171134 98132 496062
rect 99392 171134 99420 700606
rect 100772 171134 100800 700674
rect 105464 698970 105492 703520
rect 105452 698964 105504 698970
rect 105452 698906 105504 698912
rect 137848 696250 137876 703520
rect 154132 700806 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700800 154172 700806
rect 154120 700742 154172 700748
rect 137836 696244 137888 696250
rect 137836 696186 137888 696192
rect 102140 683256 102192 683262
rect 102140 683198 102192 683204
rect 98104 171106 98684 171134
rect 99392 171106 99788 171134
rect 100772 171106 100892 171134
rect 96712 170400 96764 170406
rect 96712 170342 96764 170348
rect 96620 156936 96672 156942
rect 96620 156878 96672 156884
rect 95884 155576 95936 155582
rect 95884 155518 95936 155524
rect 95608 155508 95660 155514
rect 95608 155450 95660 155456
rect 95620 153066 95648 155450
rect 95700 155440 95752 155446
rect 95700 155382 95752 155388
rect 95712 154154 95740 155382
rect 96528 154692 96580 154698
rect 96528 154634 96580 154640
rect 95700 154148 95752 154154
rect 95700 154090 95752 154096
rect 96540 154086 96568 154634
rect 96528 154080 96580 154086
rect 96528 154022 96580 154028
rect 95608 153060 95660 153066
rect 95608 153002 95660 153008
rect 96724 152674 96752 170342
rect 97632 156936 97684 156942
rect 97632 156878 97684 156884
rect 97644 152674 97672 156878
rect 98656 152674 98684 171106
rect 99760 152674 99788 171106
rect 100864 152674 100892 171106
rect 102152 152674 102180 683198
rect 103612 670744 103664 670750
rect 103612 670686 103664 670692
rect 102232 656940 102284 656946
rect 102232 656882 102284 656888
rect 102244 171134 102272 656882
rect 103624 171134 103652 670686
rect 104900 632120 104952 632126
rect 104900 632062 104952 632068
rect 104912 171134 104940 632062
rect 107660 618316 107712 618322
rect 107660 618258 107712 618264
rect 106280 605872 106332 605878
rect 106280 605814 106332 605820
rect 106292 171134 106320 605814
rect 102244 171106 103100 171134
rect 103624 171106 104204 171134
rect 104912 171106 105308 171134
rect 106292 171106 106412 171134
rect 103072 152674 103100 171106
rect 104176 152674 104204 171106
rect 105280 152674 105308 171106
rect 106384 152674 106412 171106
rect 107672 152674 107700 618258
rect 107752 579692 107804 579698
rect 107752 579634 107804 579640
rect 107764 171134 107792 579634
rect 110420 565888 110472 565894
rect 110420 565830 110472 565836
rect 109132 553444 109184 553450
rect 109132 553386 109184 553392
rect 109144 171134 109172 553386
rect 110432 171134 110460 565830
rect 111800 527196 111852 527202
rect 111800 527138 111852 527144
rect 111812 171134 111840 527138
rect 113180 514820 113232 514826
rect 113180 514762 113232 514768
rect 107764 171106 108620 171134
rect 109144 171106 109724 171134
rect 110432 171106 110828 171134
rect 111812 171106 111932 171134
rect 108592 152674 108620 171106
rect 109696 152674 109724 171106
rect 110800 152674 110828 171106
rect 111904 152674 111932 171106
rect 113192 156942 113220 514762
rect 113272 501016 113324 501022
rect 113272 500958 113324 500964
rect 113180 156936 113232 156942
rect 113180 156878 113232 156884
rect 113284 152674 113312 500958
rect 114652 474768 114704 474774
rect 114652 474710 114704 474716
rect 114664 171134 114692 474710
rect 117320 462392 117372 462398
rect 117320 462334 117372 462340
rect 115940 448588 115992 448594
rect 115940 448530 115992 448536
rect 115952 171134 115980 448530
rect 117332 171134 117360 462334
rect 120172 409896 120224 409902
rect 120172 409838 120224 409844
rect 120184 171134 120212 409838
rect 121460 371272 121512 371278
rect 121460 371214 121512 371220
rect 121472 171134 121500 371214
rect 124220 357468 124272 357474
rect 124220 357410 124272 357416
rect 122840 345092 122892 345098
rect 122840 345034 122892 345040
rect 122852 171134 122880 345034
rect 114664 171106 115244 171134
rect 115952 171106 116348 171134
rect 117332 171106 117452 171134
rect 120184 171106 120764 171134
rect 121472 171106 121868 171134
rect 122852 171106 122972 171134
rect 114192 156936 114244 156942
rect 114192 156878 114244 156884
rect 114204 152674 114232 156878
rect 115216 152674 115244 171106
rect 116320 152674 116348 171106
rect 117424 152674 117452 171106
rect 119528 162376 119580 162382
rect 119528 162318 119580 162324
rect 119540 160750 119568 162318
rect 118700 160744 118752 160750
rect 118700 160686 118752 160692
rect 119528 160744 119580 160750
rect 119528 160686 119580 160692
rect 118712 152674 118740 160686
rect 119712 158296 119764 158302
rect 119712 158238 119764 158244
rect 119724 152674 119752 158238
rect 120736 152674 120764 171106
rect 121840 152674 121868 171106
rect 122944 152674 122972 171106
rect 124232 152674 124260 357410
rect 124312 318844 124364 318850
rect 124312 318786 124364 318792
rect 124324 171134 124352 318786
rect 126980 305040 127032 305046
rect 126980 304982 127032 304988
rect 125692 292596 125744 292602
rect 125692 292538 125744 292544
rect 125704 171134 125732 292538
rect 126992 171134 127020 304982
rect 128360 266416 128412 266422
rect 128360 266358 128412 266364
rect 128372 171134 128400 266358
rect 129740 253972 129792 253978
rect 129740 253914 129792 253920
rect 124324 171106 125180 171134
rect 125704 171106 126284 171134
rect 126992 171106 127388 171134
rect 128372 171106 128492 171134
rect 125152 152674 125180 171106
rect 126256 152674 126284 171106
rect 127360 152674 127388 171106
rect 128464 152674 128492 171106
rect 129752 156942 129780 253914
rect 129832 240168 129884 240174
rect 129832 240110 129884 240116
rect 129740 156936 129792 156942
rect 129740 156878 129792 156884
rect 129844 152674 129872 240110
rect 131212 213988 131264 213994
rect 131212 213930 131264 213936
rect 131224 171134 131252 213930
rect 133880 201544 133932 201550
rect 133880 201486 133932 201492
rect 132500 187740 132552 187746
rect 132500 187682 132552 187688
rect 132512 171134 132540 187682
rect 133892 171134 133920 201486
rect 131224 171106 131804 171134
rect 132512 171106 132908 171134
rect 133892 171106 134012 171134
rect 130752 156936 130804 156942
rect 130752 156878 130804 156884
rect 130764 152674 130792 156878
rect 131776 152674 131804 171106
rect 132880 152674 132908 171106
rect 133984 152674 134012 171106
rect 135260 162920 135312 162926
rect 135260 162862 135312 162868
rect 135272 152674 135300 162862
rect 151820 162308 151872 162314
rect 151820 162250 151872 162256
rect 150716 160948 150768 160954
rect 150716 160890 150768 160896
rect 150530 158808 150586 158817
rect 150530 158743 150586 158752
rect 150438 156088 150494 156097
rect 150438 156023 150494 156032
rect 144000 155916 144052 155922
rect 144000 155858 144052 155864
rect 140780 155508 140832 155514
rect 140780 155450 140832 155456
rect 137376 155304 137428 155310
rect 137376 155246 137428 155252
rect 137192 154760 137244 154766
rect 137192 154702 137244 154708
rect 137098 154048 137154 154057
rect 137098 153983 137154 153992
rect 137112 153474 137140 153983
rect 137100 153468 137152 153474
rect 137100 153410 137152 153416
rect 137204 153134 137232 154702
rect 137284 154012 137336 154018
rect 137284 153954 137336 153960
rect 137296 153134 137324 153954
rect 137192 153128 137244 153134
rect 137192 153070 137244 153076
rect 137284 153128 137336 153134
rect 137284 153070 137336 153076
rect 137388 152674 137416 155246
rect 138020 155100 138072 155106
rect 138020 155042 138072 155048
rect 138032 154018 138060 155042
rect 140792 154630 140820 155450
rect 140964 155168 141016 155174
rect 140964 155110 141016 155116
rect 140872 154828 140924 154834
rect 140872 154770 140924 154776
rect 140780 154624 140832 154630
rect 140780 154566 140832 154572
rect 138020 154012 138072 154018
rect 138020 153954 138072 153960
rect 138480 153740 138532 153746
rect 138480 153682 138532 153688
rect 138492 152674 138520 153682
rect 140884 153202 140912 154770
rect 140872 153196 140924 153202
rect 140872 153138 140924 153144
rect 140976 152674 141004 155110
rect 142896 155032 142948 155038
rect 142896 154974 142948 154980
rect 141792 153808 141844 153814
rect 141792 153750 141844 153756
rect 141804 152674 141832 153750
rect 142908 152674 142936 154974
rect 143356 154896 143408 154902
rect 143356 154838 143408 154844
rect 143368 152969 143396 154838
rect 143448 154080 143500 154086
rect 143448 154022 143500 154028
rect 143354 152960 143410 152969
rect 143354 152895 143410 152904
rect 143460 152726 143488 154022
rect 143448 152720 143500 152726
rect 95344 152646 95772 152674
rect 96724 152646 96876 152674
rect 97644 152646 97980 152674
rect 98656 152646 99084 152674
rect 99760 152646 100188 152674
rect 100864 152646 101292 152674
rect 102152 152646 102396 152674
rect 103072 152646 103500 152674
rect 104176 152646 104604 152674
rect 105280 152646 105708 152674
rect 106384 152646 106812 152674
rect 107672 152646 107916 152674
rect 108592 152646 109020 152674
rect 109696 152646 110124 152674
rect 110800 152646 111228 152674
rect 111904 152646 112332 152674
rect 113284 152646 113436 152674
rect 114204 152646 114540 152674
rect 115216 152646 115644 152674
rect 116320 152646 116748 152674
rect 117424 152646 117852 152674
rect 118712 152646 118956 152674
rect 119724 152646 120060 152674
rect 120736 152646 121164 152674
rect 121840 152646 122268 152674
rect 122944 152646 123372 152674
rect 124232 152646 124476 152674
rect 125152 152646 125580 152674
rect 126256 152646 126684 152674
rect 127360 152646 127788 152674
rect 128464 152646 128892 152674
rect 129844 152646 129996 152674
rect 130764 152646 131100 152674
rect 131776 152646 132204 152674
rect 132880 152646 133308 152674
rect 133984 152646 134412 152674
rect 135272 152646 135516 152674
rect 137388 152646 137724 152674
rect 138492 152646 138828 152674
rect 140976 152646 141036 152674
rect 141804 152646 142140 152674
rect 142908 152646 143244 152674
rect 143448 152662 143500 152668
rect 144012 152674 144040 155858
rect 147312 155848 147364 155854
rect 147312 155790 147364 155796
rect 146300 154964 146352 154970
rect 146300 154906 146352 154912
rect 145104 154284 145156 154290
rect 145104 154226 145156 154232
rect 145116 152674 145144 154226
rect 146312 152674 146340 154906
rect 146760 154692 146812 154698
rect 146760 154634 146812 154640
rect 146772 153134 146800 154634
rect 146760 153128 146812 153134
rect 146760 153070 146812 153076
rect 147324 152674 147352 155790
rect 150452 155582 150480 156023
rect 150440 155576 150492 155582
rect 150440 155518 150492 155524
rect 150544 155310 150572 158743
rect 150532 155304 150584 155310
rect 150532 155246 150584 155252
rect 150532 154216 150584 154222
rect 150532 154158 150584 154164
rect 150440 153944 150492 153950
rect 150440 153886 150492 153892
rect 144012 152646 144348 152674
rect 145116 152646 145452 152674
rect 146312 152646 146556 152674
rect 147324 152646 147660 152674
rect 150452 152590 150480 153886
rect 150544 152658 150572 154158
rect 150532 152652 150584 152658
rect 150532 152594 150584 152600
rect 150440 152584 150492 152590
rect 95146 152552 95202 152561
rect 33046 152487 33102 152496
rect 34428 152516 34480 152522
rect 34428 152458 34480 152464
rect 35348 152516 35400 152522
rect 150440 152526 150492 152532
rect 95146 152487 95202 152496
rect 35348 152458 35400 152464
rect 34242 152416 34298 152425
rect 33948 152374 34242 152402
rect 34242 152351 34298 152360
rect 27526 152280 27582 152289
rect 27324 152238 27526 152266
rect 139596 152250 139932 152266
rect 27526 152215 27582 152224
rect 139584 152244 139932 152250
rect 139636 152238 139932 152244
rect 139584 152186 139636 152192
rect 136272 152176 136324 152182
rect 136324 152124 136620 152130
rect 136272 152118 136620 152124
rect 136284 152102 136620 152118
rect 40006 19802 40034 20060
rect 40190 19802 40218 20060
rect 40374 19802 40402 20060
rect 35808 19780 35860 19786
rect 35808 19722 35860 19728
rect 39960 19774 40034 19802
rect 40144 19774 40218 19802
rect 40328 19774 40402 19802
rect 40558 19802 40586 20060
rect 40742 19802 40770 20060
rect 40926 19802 40954 20060
rect 41110 19802 41138 20060
rect 41294 19802 41322 20060
rect 41478 19802 41506 20060
rect 40558 19774 40632 19802
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 21364 19644 21416 19650
rect 21364 19586 21416 19592
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20548 12238 20576 15574
rect 20640 14822 20668 17138
rect 21376 16318 21404 19586
rect 23388 19236 23440 19242
rect 23388 19178 23440 19184
rect 23112 17944 23164 17950
rect 23112 17886 23164 17892
rect 21364 16312 21416 16318
rect 21364 16254 21416 16260
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20916 12102 20944 15914
rect 22100 15768 22152 15774
rect 22100 15710 22152 15716
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20536 12028 20588 12034
rect 20536 11970 20588 11976
rect 20260 9240 20312 9246
rect 20260 9182 20312 9188
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 20548 9042 20576 11970
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 21100 8974 21128 14350
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21284 11354 21312 14282
rect 21364 13048 21416 13054
rect 21364 12990 21416 12996
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21376 10985 21404 12990
rect 21468 12170 21496 14554
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21362 10976 21418 10985
rect 21362 10911 21418 10920
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20640 6186 20668 8910
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20640 480 20668 3402
rect 21836 480 21864 13330
rect 22112 13161 22140 15710
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22388 14618 22416 15506
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22098 13152 22154 13161
rect 22098 13087 22154 13096
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22204 8022 22232 11562
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22756 4826 22784 11698
rect 23124 10305 23152 17886
rect 23400 15978 23428 19178
rect 23492 17678 23520 19654
rect 35820 18562 35848 19722
rect 35992 18692 36044 18698
rect 35992 18634 36044 18640
rect 36176 18692 36228 18698
rect 36176 18634 36228 18640
rect 35808 18556 35860 18562
rect 35808 18498 35860 18504
rect 33508 18488 33560 18494
rect 33508 18430 33560 18436
rect 31668 18420 31720 18426
rect 31668 18362 31720 18368
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 24872 16386 24900 17478
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25056 16574 25084 17138
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 25056 16546 25360 16574
rect 24860 16380 24912 16386
rect 24860 16322 24912 16328
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 24860 15224 24912 15230
rect 24860 15166 24912 15172
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23480 13116 23532 13122
rect 23480 13058 23532 13064
rect 23492 12034 23520 13058
rect 23480 12028 23532 12034
rect 23480 11970 23532 11976
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23110 10296 23166 10305
rect 23110 10231 23166 10240
rect 23492 7614 23520 10610
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23480 7608 23532 7614
rect 23480 7550 23532 7556
rect 23584 7138 23612 10542
rect 23676 9586 23704 13466
rect 24872 13122 24900 15166
rect 24860 13116 24912 13122
rect 24860 13058 24912 13064
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23768 9489 23796 12106
rect 24872 10878 24900 12174
rect 24860 10872 24912 10878
rect 24860 10814 24912 10820
rect 23754 9480 23810 9489
rect 23754 9415 23810 9424
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 23572 7132 23624 7138
rect 23572 7074 23624 7080
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 23032 480 23060 6394
rect 24228 480 24256 7754
rect 25332 480 25360 16546
rect 26252 16454 26280 17070
rect 27620 16856 27672 16862
rect 27620 16798 27672 16804
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 27632 13870 27660 16798
rect 27724 16574 27752 17478
rect 27724 16546 28488 16574
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 11630
rect 26332 9308 26384 9314
rect 26332 9250 26384 9256
rect 26344 6254 26372 9250
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 27712 4956 27764 4962
rect 27712 4898 27764 4904
rect 27724 480 27752 4898
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 29104 7886 29132 10678
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 30116 480 30144 10610
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 14350
rect 31680 13462 31708 18362
rect 33520 13530 33548 18430
rect 33692 15836 33744 15842
rect 33692 15778 33744 15784
rect 33508 13524 33560 13530
rect 33508 13466 33560 13472
rect 31668 13456 31720 13462
rect 31668 13398 31720 13404
rect 33704 13122 33732 15778
rect 33876 13864 33928 13870
rect 33876 13806 33928 13812
rect 33140 13116 33192 13122
rect 33140 13058 33192 13064
rect 33692 13116 33744 13122
rect 33692 13058 33744 13064
rect 33152 10742 33180 13058
rect 33140 10736 33192 10742
rect 33140 10678 33192 10684
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 32416 480 32444 3538
rect 33152 2786 33180 6258
rect 33888 6225 33916 13806
rect 36004 11665 36032 18634
rect 36188 17610 36216 18634
rect 36176 17604 36228 17610
rect 36176 17546 36228 17552
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 35990 11656 36046 11665
rect 35990 11591 36046 11600
rect 35900 7676 35952 7682
rect 35900 7618 35952 7624
rect 35912 6905 35940 7618
rect 35898 6896 35954 6905
rect 35898 6831 35954 6840
rect 33874 6216 33930 6225
rect 33874 6151 33930 6160
rect 36556 3874 36584 17206
rect 39304 16720 39356 16726
rect 39304 16662 39356 16668
rect 37188 13524 37240 13530
rect 37188 13466 37240 13472
rect 36820 13456 36872 13462
rect 36820 13398 36872 13404
rect 36832 7682 36860 13398
rect 37200 7954 37228 13466
rect 37188 7948 37240 7954
rect 37188 7890 37240 7896
rect 36820 7676 36872 7682
rect 36820 7618 36872 7624
rect 33600 3868 33652 3874
rect 33600 3810 33652 3816
rect 36544 3868 36596 3874
rect 36544 3810 36596 3816
rect 33140 2780 33192 2786
rect 33140 2722 33192 2728
rect 33612 480 33640 3810
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34808 480 34836 3742
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 35992 3324 36044 3330
rect 35992 3266 36044 3272
rect 36004 480 36032 3266
rect 37188 2984 37240 2990
rect 37188 2926 37240 2932
rect 37200 480 37228 2926
rect 38396 480 38424 3470
rect 39316 3330 39344 16662
rect 39960 16046 39988 19774
rect 40040 17604 40092 17610
rect 40040 17546 40092 17552
rect 39948 16040 40000 16046
rect 39948 15982 40000 15988
rect 40052 13326 40080 17546
rect 40144 15910 40172 19774
rect 40328 16402 40356 19774
rect 40236 16374 40356 16402
rect 40132 15904 40184 15910
rect 40132 15846 40184 15852
rect 40236 14482 40264 16374
rect 40604 14498 40632 19774
rect 40224 14476 40276 14482
rect 40224 14418 40276 14424
rect 40316 14476 40368 14482
rect 40316 14418 40368 14424
rect 40512 14470 40632 14498
rect 40696 19774 40770 19802
rect 40880 19774 40954 19802
rect 41064 19774 41138 19802
rect 41248 19774 41322 19802
rect 41432 19774 41506 19802
rect 41662 19802 41690 20060
rect 41846 19802 41874 20060
rect 42030 19938 42058 20060
rect 42030 19910 42104 19938
rect 41662 19774 41736 19802
rect 40696 14482 40724 19774
rect 40776 17944 40828 17950
rect 40776 17886 40828 17892
rect 40684 14476 40736 14482
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 40328 6390 40356 14418
rect 40512 7750 40540 14470
rect 40684 14418 40736 14424
rect 40592 13252 40644 13258
rect 40592 13194 40644 13200
rect 40604 10606 40632 13194
rect 40684 11960 40736 11966
rect 40684 11902 40736 11908
rect 40592 10600 40644 10606
rect 40592 10542 40644 10548
rect 40500 7744 40552 7750
rect 40500 7686 40552 7692
rect 40316 6384 40368 6390
rect 40316 6326 40368 6332
rect 40696 3670 40724 11902
rect 40788 9178 40816 17886
rect 40880 16998 40908 19774
rect 40868 16992 40920 16998
rect 40868 16934 40920 16940
rect 41064 16114 41092 19774
rect 41052 16108 41104 16114
rect 41052 16050 41104 16056
rect 41248 11898 41276 19774
rect 41432 17338 41460 19774
rect 41604 18420 41656 18426
rect 41604 18362 41656 18368
rect 41420 17332 41472 17338
rect 41420 17274 41472 17280
rect 41616 16182 41644 18362
rect 41604 16176 41656 16182
rect 41604 16118 41656 16124
rect 41236 11892 41288 11898
rect 41236 11834 41288 11840
rect 40776 9172 40828 9178
rect 40776 9114 40828 9120
rect 41708 4894 41736 19774
rect 41800 19774 41874 19802
rect 41800 18426 41828 19774
rect 41788 18420 41840 18426
rect 41788 18362 41840 18368
rect 42076 17950 42104 19910
rect 42214 19802 42242 20060
rect 42398 19802 42426 20060
rect 42582 19802 42610 20060
rect 42766 19802 42794 20060
rect 42950 19938 42978 20060
rect 42950 19910 43024 19938
rect 42168 19774 42242 19802
rect 42352 19774 42426 19802
rect 42536 19774 42610 19802
rect 42720 19774 42794 19802
rect 42064 17944 42116 17950
rect 42064 17886 42116 17892
rect 42168 17762 42196 19774
rect 41800 17734 42196 17762
rect 41800 10538 41828 17734
rect 42352 17406 42380 19774
rect 42340 17400 42392 17406
rect 42340 17342 42392 17348
rect 42064 17128 42116 17134
rect 42064 17070 42116 17076
rect 41788 10532 41840 10538
rect 41788 10474 41840 10480
rect 41696 4888 41748 4894
rect 41696 4830 41748 4836
rect 40684 3664 40736 3670
rect 40684 3606 40736 3612
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 39304 3324 39356 3330
rect 39304 3266 39356 3272
rect 39580 3188 39632 3194
rect 39580 3130 39632 3136
rect 39592 480 39620 3130
rect 40696 480 40724 3402
rect 41892 480 41920 3538
rect 42076 3194 42104 17070
rect 42156 17060 42208 17066
rect 42156 17002 42208 17008
rect 42168 3534 42196 17002
rect 42248 15224 42300 15230
rect 42248 15166 42300 15172
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42260 3398 42288 15166
rect 42536 14550 42564 19774
rect 42720 17610 42748 19774
rect 42892 18420 42944 18426
rect 42892 18362 42944 18368
rect 42708 17604 42760 17610
rect 42708 17546 42760 17552
rect 42904 15230 42932 18362
rect 42996 17474 43024 19910
rect 43134 19802 43162 20060
rect 43088 19774 43162 19802
rect 43318 19802 43346 20060
rect 43502 19802 43530 20060
rect 43686 19802 43714 20060
rect 43870 19802 43898 20060
rect 44054 19802 44082 20060
rect 43318 19774 43392 19802
rect 43088 18426 43116 19774
rect 43076 18420 43128 18426
rect 43076 18362 43128 18368
rect 43364 18170 43392 19774
rect 43168 18148 43220 18154
rect 43168 18090 43220 18096
rect 43272 18142 43392 18170
rect 43456 19774 43530 19802
rect 43640 19774 43714 19802
rect 43824 19774 43898 19802
rect 44008 19774 44082 19802
rect 44238 19802 44266 20060
rect 44422 19938 44450 20060
rect 44422 19910 44496 19938
rect 44238 19774 44404 19802
rect 43076 18080 43128 18086
rect 43076 18022 43128 18028
rect 42984 17468 43036 17474
rect 42984 17410 43036 17416
rect 42892 15224 42944 15230
rect 42892 15166 42944 15172
rect 42524 14544 42576 14550
rect 42524 14486 42576 14492
rect 42800 10736 42852 10742
rect 42800 10678 42852 10684
rect 42812 7750 42840 10678
rect 42800 7744 42852 7750
rect 42800 7686 42852 7692
rect 43088 6458 43116 18022
rect 43180 7818 43208 18090
rect 43272 13394 43300 18142
rect 43456 18086 43484 19774
rect 43640 18154 43668 19774
rect 43628 18148 43680 18154
rect 43628 18090 43680 18096
rect 43444 18080 43496 18086
rect 43444 18022 43496 18028
rect 43352 17604 43404 17610
rect 43352 17546 43404 17552
rect 43364 16250 43392 17546
rect 43444 17332 43496 17338
rect 43444 17274 43496 17280
rect 43352 16244 43404 16250
rect 43352 16186 43404 16192
rect 43260 13388 43312 13394
rect 43260 13330 43312 13336
rect 43168 7812 43220 7818
rect 43168 7754 43220 7760
rect 43076 6452 43128 6458
rect 43076 6394 43128 6400
rect 43076 3868 43128 3874
rect 43076 3810 43128 3816
rect 42248 3392 42300 3398
rect 42248 3334 42300 3340
rect 42064 3188 42116 3194
rect 42064 3130 42116 3136
rect 43088 480 43116 3810
rect 43456 3738 43484 17274
rect 43824 17202 43852 19774
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 43536 16856 43588 16862
rect 43536 16798 43588 16804
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 43548 2990 43576 16798
rect 43628 16788 43680 16794
rect 43628 16730 43680 16736
rect 43640 3466 43668 16730
rect 44008 11694 44036 19774
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 44192 16574 44220 16934
rect 44192 16546 44312 16574
rect 43996 11688 44048 11694
rect 43996 11630 44048 11636
rect 43628 3460 43680 3466
rect 43628 3402 43680 3408
rect 43536 2984 43588 2990
rect 43536 2926 43588 2932
rect 44284 480 44312 16546
rect 44376 4962 44404 19774
rect 44468 17542 44496 19910
rect 44606 19802 44634 20060
rect 44790 19802 44818 20060
rect 44974 19802 45002 20060
rect 45158 19802 45186 20060
rect 45342 19802 45370 20060
rect 45526 19802 45554 20060
rect 45710 19802 45738 20060
rect 45894 19802 45922 20060
rect 46078 19802 46106 20060
rect 46262 19802 46290 20060
rect 46446 19802 46474 20060
rect 46630 19802 46658 20060
rect 46814 19802 46842 20060
rect 44560 19774 44634 19802
rect 44744 19774 44818 19802
rect 44928 19774 45002 19802
rect 45112 19774 45186 19802
rect 45296 19774 45370 19802
rect 45480 19774 45554 19802
rect 45664 19774 45738 19802
rect 45848 19774 45922 19802
rect 46032 19774 46106 19802
rect 46216 19774 46290 19802
rect 46400 19774 46474 19802
rect 46584 19774 46658 19802
rect 46768 19774 46842 19802
rect 46998 19802 47026 20060
rect 47182 19802 47210 20060
rect 47366 19802 47394 20060
rect 47550 19802 47578 20060
rect 46998 19774 47072 19802
rect 44456 17536 44508 17542
rect 44456 17478 44508 17484
rect 44560 10674 44588 19774
rect 44744 14414 44772 19774
rect 44928 17338 44956 19774
rect 44916 17332 44968 17338
rect 44916 17274 44968 17280
rect 45112 17270 45140 19774
rect 45100 17264 45152 17270
rect 45100 17206 45152 17212
rect 44824 16652 44876 16658
rect 44824 16594 44876 16600
rect 44732 14408 44784 14414
rect 44732 14350 44784 14356
rect 44548 10668 44600 10674
rect 44548 10610 44600 10616
rect 44364 4956 44416 4962
rect 44364 4898 44416 4904
rect 44836 3602 44864 16594
rect 45296 3806 45324 19774
rect 45480 16726 45508 19774
rect 45560 17944 45612 17950
rect 45560 17886 45612 17892
rect 45468 16720 45520 16726
rect 45468 16662 45520 16668
rect 45572 6914 45600 17886
rect 45664 16862 45692 19774
rect 45744 17400 45796 17406
rect 45744 17342 45796 17348
rect 45652 16856 45704 16862
rect 45652 16798 45704 16804
rect 45756 15502 45784 17342
rect 45848 17066 45876 19774
rect 46032 17134 46060 19774
rect 46020 17128 46072 17134
rect 46020 17070 46072 17076
rect 45836 17060 45888 17066
rect 45836 17002 45888 17008
rect 46216 16794 46244 19774
rect 46204 16788 46256 16794
rect 46204 16730 46256 16736
rect 46400 16658 46428 19774
rect 46388 16652 46440 16658
rect 46388 16594 46440 16600
rect 45744 15496 45796 15502
rect 45744 15438 45796 15444
rect 45572 6886 46520 6914
rect 45284 3800 45336 3806
rect 45284 3742 45336 3748
rect 44824 3596 44876 3602
rect 44824 3538 44876 3544
rect 46492 3482 46520 6886
rect 46584 3874 46612 19774
rect 46768 16998 46796 19774
rect 46756 16992 46808 16998
rect 46756 16934 46808 16940
rect 46572 3868 46624 3874
rect 46572 3810 46624 3816
rect 45468 3460 45520 3466
rect 46492 3454 46704 3482
rect 47044 3466 47072 19774
rect 47136 19774 47210 19802
rect 47320 19774 47394 19802
rect 47504 19774 47578 19802
rect 47734 19802 47762 20060
rect 47918 19802 47946 20060
rect 48102 19802 48130 20060
rect 48286 19802 48314 20060
rect 47734 19774 47808 19802
rect 47918 19774 47992 19802
rect 48102 19774 48176 19802
rect 47136 17950 47164 19774
rect 47124 17944 47176 17950
rect 47124 17886 47176 17892
rect 47320 16574 47348 19774
rect 47320 16546 47440 16574
rect 47308 16176 47360 16182
rect 47308 16118 47360 16124
rect 47320 14618 47348 16118
rect 47308 14612 47360 14618
rect 47308 14554 47360 14560
rect 45468 3402 45520 3408
rect 45480 480 45508 3402
rect 46676 480 46704 3454
rect 47032 3460 47084 3466
rect 47032 3402 47084 3408
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47504 3466 47532 19774
rect 47780 17202 47808 19774
rect 47964 17338 47992 19774
rect 47952 17332 48004 17338
rect 47952 17274 48004 17280
rect 47768 17196 47820 17202
rect 47768 17138 47820 17144
rect 48148 17066 48176 19774
rect 48240 19774 48314 19802
rect 48470 19802 48498 20060
rect 48654 19802 48682 20060
rect 48838 19802 48866 20060
rect 49022 19802 49050 20060
rect 49206 19802 49234 20060
rect 49390 19802 49418 20060
rect 49574 19802 49602 20060
rect 48470 19774 48544 19802
rect 48654 19774 48728 19802
rect 48838 19774 48912 19802
rect 48240 17270 48268 19774
rect 48516 17950 48544 19774
rect 48504 17944 48556 17950
rect 48504 17886 48556 17892
rect 48228 17264 48280 17270
rect 48228 17206 48280 17212
rect 48136 17060 48188 17066
rect 48136 17002 48188 17008
rect 48700 16998 48728 19774
rect 48884 17134 48912 19774
rect 48976 19774 49050 19802
rect 49160 19774 49234 19802
rect 49344 19774 49418 19802
rect 49528 19774 49602 19802
rect 49758 19802 49786 20060
rect 49942 19802 49970 20060
rect 50126 19802 50154 20060
rect 49758 19774 49832 19802
rect 48872 17128 48924 17134
rect 48872 17070 48924 17076
rect 48688 16992 48740 16998
rect 48688 16934 48740 16940
rect 48976 3738 49004 19774
rect 48964 3732 49016 3738
rect 48964 3674 49016 3680
rect 47492 3460 47544 3466
rect 47492 3402 47544 3408
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48976 480 49004 3402
rect 49160 3330 49188 19774
rect 49344 3670 49372 19774
rect 49528 3806 49556 19774
rect 49804 17202 49832 19774
rect 49896 19774 49970 19802
rect 50080 19774 50154 19802
rect 50310 19802 50338 20060
rect 50494 19802 50522 20060
rect 50678 19802 50706 20060
rect 50862 19802 50890 20060
rect 51046 19802 51074 20060
rect 50310 19774 50384 19802
rect 49700 17196 49752 17202
rect 49700 17138 49752 17144
rect 49792 17196 49844 17202
rect 49792 17138 49844 17144
rect 49712 6914 49740 17138
rect 49896 8906 49924 19774
rect 50080 15774 50108 19774
rect 50356 17474 50384 19774
rect 50448 19774 50522 19802
rect 50632 19774 50706 19802
rect 50816 19774 50890 19802
rect 51000 19774 51074 19802
rect 51230 19802 51258 20060
rect 51414 19802 51442 20060
rect 51598 19802 51626 20060
rect 51782 19802 51810 20060
rect 51966 19802 51994 20060
rect 51230 19774 51304 19802
rect 51414 19774 51488 19802
rect 50344 17468 50396 17474
rect 50344 17410 50396 17416
rect 50344 17332 50396 17338
rect 50344 17274 50396 17280
rect 50068 15768 50120 15774
rect 50068 15710 50120 15716
rect 49884 8900 49936 8906
rect 49884 8842 49936 8848
rect 49712 6886 50200 6914
rect 49516 3800 49568 3806
rect 49516 3742 49568 3748
rect 49332 3664 49384 3670
rect 49332 3606 49384 3612
rect 49148 3324 49200 3330
rect 49148 3266 49200 3272
rect 50172 480 50200 6886
rect 50356 3466 50384 17274
rect 50448 11898 50476 19774
rect 50528 17060 50580 17066
rect 50528 17002 50580 17008
rect 50436 11892 50488 11898
rect 50436 11834 50488 11840
rect 50540 3602 50568 17002
rect 50632 6594 50660 19774
rect 50712 17944 50764 17950
rect 50712 17886 50764 17892
rect 50620 6588 50672 6594
rect 50620 6530 50672 6536
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50344 3460 50396 3466
rect 50344 3402 50396 3408
rect 50724 3398 50752 17886
rect 50816 14210 50844 19774
rect 50804 14204 50856 14210
rect 50804 14146 50856 14152
rect 51000 13394 51028 19774
rect 51276 17610 51304 19774
rect 51264 17604 51316 17610
rect 51264 17546 51316 17552
rect 51460 16862 51488 19774
rect 51552 19774 51626 19802
rect 51736 19774 51810 19802
rect 51920 19774 51994 19802
rect 52150 19802 52178 20060
rect 52334 19802 52362 20060
rect 52150 19774 52224 19802
rect 51448 16856 51500 16862
rect 51448 16798 51500 16804
rect 50988 13388 51040 13394
rect 50988 13330 51040 13336
rect 51552 13326 51580 19774
rect 51540 13320 51592 13326
rect 51540 13262 51592 13268
rect 51736 10742 51764 19774
rect 51816 17468 51868 17474
rect 51816 17410 51868 17416
rect 51724 10736 51776 10742
rect 51724 10678 51776 10684
rect 51828 5166 51856 17410
rect 51816 5160 51868 5166
rect 51816 5102 51868 5108
rect 51920 5030 51948 19774
rect 52196 17950 52224 19774
rect 52288 19774 52362 19802
rect 52518 19802 52546 20060
rect 52702 19802 52730 20060
rect 52886 19802 52914 20060
rect 53070 19802 53098 20060
rect 53254 19802 53282 20060
rect 53438 19802 53466 20060
rect 52518 19774 52592 19802
rect 52702 19774 52776 19802
rect 52184 17944 52236 17950
rect 52184 17886 52236 17892
rect 52288 6458 52316 19774
rect 52460 17944 52512 17950
rect 52460 17886 52512 17892
rect 52472 10198 52500 17886
rect 52564 16794 52592 19774
rect 52748 17474 52776 19774
rect 52840 19774 52914 19802
rect 53024 19774 53098 19802
rect 53208 19774 53282 19802
rect 53392 19774 53466 19802
rect 53622 19802 53650 20060
rect 53806 19802 53834 20060
rect 53990 19802 54018 20060
rect 54174 19802 54202 20060
rect 54358 19802 54386 20060
rect 54542 19802 54570 20060
rect 54726 19802 54754 20060
rect 53622 19774 53696 19802
rect 52736 17468 52788 17474
rect 52736 17410 52788 17416
rect 52736 17264 52788 17270
rect 52736 17206 52788 17212
rect 52552 16788 52604 16794
rect 52552 16730 52604 16736
rect 52460 10192 52512 10198
rect 52460 10134 52512 10140
rect 52748 6914 52776 17206
rect 52840 9382 52868 19774
rect 52828 9376 52880 9382
rect 52828 9318 52880 9324
rect 52748 6886 52960 6914
rect 52276 6452 52328 6458
rect 52276 6394 52328 6400
rect 51908 5024 51960 5030
rect 51908 4966 51960 4972
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 50712 3392 50764 3398
rect 50712 3334 50764 3340
rect 51368 480 51396 3402
rect 52564 480 52592 3538
rect 52932 490 52960 6886
rect 53024 4962 53052 19774
rect 53104 17604 53156 17610
rect 53104 17546 53156 17552
rect 53116 6526 53144 17546
rect 53208 15706 53236 19774
rect 53196 15700 53248 15706
rect 53196 15642 53248 15648
rect 53104 6520 53156 6526
rect 53104 6462 53156 6468
rect 53392 6390 53420 19774
rect 53668 17066 53696 19774
rect 53760 19774 53834 19802
rect 53944 19774 54018 19802
rect 54128 19774 54202 19802
rect 54312 19774 54386 19802
rect 54496 19774 54570 19802
rect 54680 19774 54754 19802
rect 54910 19802 54938 20060
rect 55094 19802 55122 20060
rect 55278 19802 55306 20060
rect 55462 19802 55490 20060
rect 55646 19802 55674 20060
rect 55830 19802 55858 20060
rect 56014 19802 56042 20060
rect 56198 19802 56226 20060
rect 56382 19802 56410 20060
rect 56566 19802 56594 20060
rect 56750 19802 56778 20060
rect 56934 19802 56962 20060
rect 57118 19802 57146 20060
rect 57302 19802 57330 20060
rect 54910 19774 54984 19802
rect 53656 17060 53708 17066
rect 53656 17002 53708 17008
rect 53760 13530 53788 19774
rect 53944 16114 53972 19774
rect 53932 16108 53984 16114
rect 53932 16050 53984 16056
rect 54128 14550 54156 19774
rect 54116 14544 54168 14550
rect 54116 14486 54168 14492
rect 53748 13524 53800 13530
rect 53748 13466 53800 13472
rect 54312 7818 54340 19774
rect 54496 10062 54524 19774
rect 54576 17128 54628 17134
rect 54576 17070 54628 17076
rect 54484 10056 54536 10062
rect 54484 9998 54536 10004
rect 54300 7812 54352 7818
rect 54300 7754 54352 7760
rect 53380 6384 53432 6390
rect 53380 6326 53432 6332
rect 53012 4956 53064 4962
rect 53012 4898 53064 4904
rect 54588 4146 54616 17070
rect 54680 13258 54708 19774
rect 54956 17338 54984 19774
rect 55048 19774 55122 19802
rect 55232 19774 55306 19802
rect 55416 19774 55490 19802
rect 55600 19774 55674 19802
rect 55784 19774 55858 19802
rect 55968 19774 56042 19802
rect 56152 19774 56226 19802
rect 56336 19774 56410 19802
rect 56520 19774 56594 19802
rect 56704 19774 56778 19802
rect 56888 19774 56962 19802
rect 57072 19774 57146 19802
rect 57256 19774 57330 19802
rect 57486 19802 57514 20060
rect 57670 19802 57698 20060
rect 57854 19802 57882 20060
rect 58038 19802 58066 20060
rect 58222 19802 58250 20060
rect 58406 19802 58434 20060
rect 58590 19802 58618 20060
rect 58774 19802 58802 20060
rect 58958 19802 58986 20060
rect 57486 19774 57560 19802
rect 54944 17332 54996 17338
rect 54944 17274 54996 17280
rect 54944 17060 54996 17066
rect 54944 17002 54996 17008
rect 54760 16992 54812 16998
rect 54760 16934 54812 16940
rect 54668 13252 54720 13258
rect 54668 13194 54720 13200
rect 54576 4140 54628 4146
rect 54576 4082 54628 4088
rect 54772 3466 54800 16934
rect 54956 4894 54984 17002
rect 55048 9178 55076 19774
rect 55232 14482 55260 19774
rect 55416 16046 55444 19774
rect 55600 16250 55628 19774
rect 55588 16244 55640 16250
rect 55588 16186 55640 16192
rect 55404 16040 55456 16046
rect 55404 15982 55456 15988
rect 55220 14476 55272 14482
rect 55220 14418 55272 14424
rect 55784 10538 55812 19774
rect 55864 16788 55916 16794
rect 55864 16730 55916 16736
rect 55772 10532 55824 10538
rect 55772 10474 55824 10480
rect 55036 9172 55088 9178
rect 55036 9114 55088 9120
rect 55876 5098 55904 16730
rect 55968 11966 55996 19774
rect 56048 16856 56100 16862
rect 56048 16798 56100 16804
rect 55956 11960 56008 11966
rect 55956 11902 56008 11908
rect 55864 5092 55916 5098
rect 55864 5034 55916 5040
rect 54944 4888 54996 4894
rect 54944 4830 54996 4836
rect 56060 4758 56088 16798
rect 56152 10674 56180 19774
rect 56336 15842 56364 19774
rect 56520 17134 56548 19774
rect 56508 17128 56560 17134
rect 56508 17070 56560 17076
rect 56324 15836 56376 15842
rect 56324 15778 56376 15784
rect 56140 10668 56192 10674
rect 56140 10610 56192 10616
rect 56600 9240 56652 9246
rect 56600 9182 56652 9188
rect 56612 6866 56640 9182
rect 56704 8838 56732 19774
rect 56888 11694 56916 19774
rect 57072 14618 57100 19774
rect 57060 14612 57112 14618
rect 57060 14554 57112 14560
rect 56876 11688 56928 11694
rect 56876 11630 56928 11636
rect 56692 8832 56744 8838
rect 56692 8774 56744 8780
rect 56600 6860 56652 6866
rect 56600 6802 56652 6808
rect 57256 6322 57284 19774
rect 57532 17610 57560 19774
rect 57624 19774 57698 19802
rect 57808 19774 57882 19802
rect 57992 19774 58066 19802
rect 58176 19774 58250 19802
rect 58360 19774 58434 19802
rect 58544 19774 58618 19802
rect 58728 19774 58802 19802
rect 58912 19774 58986 19802
rect 59142 19802 59170 20060
rect 59326 19802 59354 20060
rect 59510 19802 59538 20060
rect 59694 19802 59722 20060
rect 59878 19802 59906 20060
rect 59142 19774 59216 19802
rect 57520 17604 57572 17610
rect 57520 17546 57572 17552
rect 57624 15910 57652 19774
rect 57612 15904 57664 15910
rect 57612 15846 57664 15852
rect 57336 13524 57388 13530
rect 57336 13466 57388 13472
rect 57244 6316 57296 6322
rect 57244 6258 57296 6264
rect 56508 4820 56560 4826
rect 56508 4762 56560 4768
rect 56048 4752 56100 4758
rect 56048 4694 56100 4700
rect 54760 3460 54812 3466
rect 54760 3402 54812 3408
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 54944 3392 54996 3398
rect 54944 3334 54996 3340
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 52932 462 53328 490
rect 54956 480 54984 3334
rect 56060 480 56088 3402
rect 56520 2417 56548 4762
rect 57244 4140 57296 4146
rect 57244 4082 57296 4088
rect 56506 2408 56562 2417
rect 56506 2343 56562 2352
rect 57256 480 57284 4082
rect 57348 3738 57376 13466
rect 57808 11626 57836 19774
rect 57796 11620 57848 11626
rect 57796 11562 57848 11568
rect 57888 10464 57940 10470
rect 57888 10406 57940 10412
rect 57900 7206 57928 10406
rect 57992 7342 58020 19774
rect 58176 14958 58204 19774
rect 58164 14952 58216 14958
rect 58164 14894 58216 14900
rect 58360 11558 58388 19774
rect 58544 12918 58572 19774
rect 58728 14142 58756 19774
rect 58716 14136 58768 14142
rect 58716 14078 58768 14084
rect 58532 12912 58584 12918
rect 58532 12854 58584 12860
rect 58348 11552 58400 11558
rect 58348 11494 58400 11500
rect 57980 7336 58032 7342
rect 57980 7278 58032 7284
rect 57888 7200 57940 7206
rect 57888 7142 57940 7148
rect 57336 3732 57388 3738
rect 57336 3674 57388 3680
rect 58440 3664 58492 3670
rect 58440 3606 58492 3612
rect 58452 480 58480 3606
rect 58912 2514 58940 19774
rect 59188 16574 59216 19774
rect 59096 16546 59216 16574
rect 59280 19774 59354 19802
rect 59464 19774 59538 19802
rect 59648 19774 59722 19802
rect 59832 19774 59906 19802
rect 60062 19802 60090 20060
rect 60246 19802 60274 20060
rect 60430 19802 60458 20060
rect 60614 19802 60642 20060
rect 60062 19774 60136 19802
rect 59096 12782 59124 16546
rect 59176 15972 59228 15978
rect 59176 15914 59228 15920
rect 59188 13705 59216 15914
rect 59174 13696 59230 13705
rect 59174 13631 59230 13640
rect 59084 12776 59136 12782
rect 59084 12718 59136 12724
rect 59280 6914 59308 19774
rect 59188 6886 59308 6914
rect 59188 4078 59216 6886
rect 59268 6180 59320 6186
rect 59268 6122 59320 6128
rect 59280 4554 59308 6122
rect 59464 5302 59492 19774
rect 59648 5574 59676 19774
rect 59832 10946 59860 19774
rect 60108 19242 60136 19774
rect 60200 19774 60274 19802
rect 60384 19774 60458 19802
rect 60568 19774 60642 19802
rect 60798 19802 60826 20060
rect 60982 19802 61010 20060
rect 60798 19774 60872 19802
rect 60096 19236 60148 19242
rect 60096 19178 60148 19184
rect 60004 17264 60056 17270
rect 60004 17206 60056 17212
rect 59820 10940 59872 10946
rect 59820 10882 59872 10888
rect 59912 10396 59964 10402
rect 59912 10338 59964 10344
rect 59924 8498 59952 10338
rect 59912 8492 59964 8498
rect 59912 8434 59964 8440
rect 59636 5568 59688 5574
rect 59636 5510 59688 5516
rect 59452 5296 59504 5302
rect 59452 5238 59504 5244
rect 59268 4548 59320 4554
rect 59268 4490 59320 4496
rect 59176 4072 59228 4078
rect 59176 4014 59228 4020
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 58900 2508 58952 2514
rect 58900 2450 58952 2456
rect 59648 480 59676 3334
rect 60016 3262 60044 17206
rect 60200 15230 60228 19774
rect 60188 15224 60240 15230
rect 60188 15166 60240 15172
rect 60096 14612 60148 14618
rect 60096 14554 60148 14560
rect 60108 3466 60136 14554
rect 60384 14414 60412 19774
rect 60372 14408 60424 14414
rect 60372 14350 60424 14356
rect 60568 4570 60596 19774
rect 60648 17944 60700 17950
rect 60648 17886 60700 17892
rect 60660 14686 60688 17886
rect 60844 17202 60872 19774
rect 60936 19774 61010 19802
rect 61166 19802 61194 20060
rect 61350 19802 61378 20060
rect 61534 19802 61562 20060
rect 61166 19774 61240 19802
rect 60832 17196 60884 17202
rect 60832 17138 60884 17144
rect 60648 14680 60700 14686
rect 60648 14622 60700 14628
rect 60936 10266 60964 19774
rect 61212 18902 61240 19774
rect 61304 19774 61378 19802
rect 61488 19774 61562 19802
rect 61718 19802 61746 20060
rect 61902 19938 61930 20060
rect 61856 19910 61930 19938
rect 61718 19774 61792 19802
rect 61200 18896 61252 18902
rect 61200 18838 61252 18844
rect 61304 14346 61332 19774
rect 61384 17332 61436 17338
rect 61384 17274 61436 17280
rect 61292 14340 61344 14346
rect 61292 14282 61344 14288
rect 60924 10260 60976 10266
rect 60924 10202 60976 10208
rect 60924 5296 60976 5302
rect 60924 5238 60976 5244
rect 60568 4542 60780 4570
rect 60096 3460 60148 3466
rect 60096 3402 60148 3408
rect 60004 3256 60056 3262
rect 60004 3198 60056 3204
rect 60752 2174 60780 4542
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 60740 2168 60792 2174
rect 60740 2110 60792 2116
rect 60844 480 60872 3538
rect 60936 950 60964 5238
rect 61396 3670 61424 17274
rect 61488 10402 61516 19774
rect 61660 16720 61712 16726
rect 61660 16662 61712 16668
rect 61568 15700 61620 15706
rect 61568 15642 61620 15648
rect 61476 10396 61528 10402
rect 61476 10338 61528 10344
rect 61580 3874 61608 15642
rect 61672 14754 61700 16662
rect 61764 16658 61792 19774
rect 61856 17338 61884 19910
rect 62086 19802 62114 20060
rect 61948 19774 62114 19802
rect 62270 19802 62298 20060
rect 62454 19802 62482 20060
rect 62638 19802 62666 20060
rect 62822 19802 62850 20060
rect 63006 19802 63034 20060
rect 63190 19802 63218 20060
rect 63374 19802 63402 20060
rect 63558 19802 63586 20060
rect 62270 19774 62344 19802
rect 61844 17332 61896 17338
rect 61844 17274 61896 17280
rect 61752 16652 61804 16658
rect 61752 16594 61804 16600
rect 61844 15224 61896 15230
rect 61844 15166 61896 15172
rect 61660 14748 61712 14754
rect 61660 14690 61712 14696
rect 61660 10940 61712 10946
rect 61660 10882 61712 10888
rect 61672 7478 61700 10882
rect 61856 7546 61884 15166
rect 61948 10470 61976 19774
rect 62316 19106 62344 19774
rect 62408 19774 62482 19802
rect 62592 19774 62666 19802
rect 62776 19774 62850 19802
rect 62960 19774 63034 19802
rect 63144 19774 63218 19802
rect 63328 19774 63402 19802
rect 63512 19774 63586 19802
rect 63742 19802 63770 20060
rect 63926 19802 63954 20060
rect 64110 19802 64138 20060
rect 64294 19802 64322 20060
rect 64478 19802 64506 20060
rect 64662 19802 64690 20060
rect 64846 19802 64874 20060
rect 65030 19802 65058 20060
rect 65214 19802 65242 20060
rect 65398 19802 65426 20060
rect 65582 19802 65610 20060
rect 63742 19774 63816 19802
rect 63926 19774 64000 19802
rect 64110 19774 64184 19802
rect 64294 19774 64368 19802
rect 64478 19774 64552 19802
rect 64662 19774 64736 19802
rect 62304 19100 62356 19106
rect 62304 19042 62356 19048
rect 62028 17604 62080 17610
rect 62028 17546 62080 17552
rect 62040 15774 62068 17546
rect 62028 15768 62080 15774
rect 62028 15710 62080 15716
rect 61936 10464 61988 10470
rect 61936 10406 61988 10412
rect 61844 7540 61896 7546
rect 61844 7482 61896 7488
rect 61660 7472 61712 7478
rect 61660 7414 61712 7420
rect 62408 6050 62436 19774
rect 62396 6044 62448 6050
rect 62396 5986 62448 5992
rect 62592 4486 62620 19774
rect 62776 14890 62804 19774
rect 62960 17542 62988 19774
rect 62948 17536 63000 17542
rect 62948 17478 63000 17484
rect 62764 14884 62816 14890
rect 62764 14826 62816 14832
rect 63144 10878 63172 19774
rect 63328 17950 63356 19774
rect 63408 19372 63460 19378
rect 63408 19314 63460 19320
rect 63420 18222 63448 19314
rect 63408 18216 63460 18222
rect 63408 18158 63460 18164
rect 63316 17944 63368 17950
rect 63316 17886 63368 17892
rect 63132 10872 63184 10878
rect 63132 10814 63184 10820
rect 62580 4480 62632 4486
rect 62580 4422 62632 4428
rect 61568 3868 61620 3874
rect 61568 3810 61620 3816
rect 62028 3800 62080 3806
rect 62028 3742 62080 3748
rect 61384 3664 61436 3670
rect 61384 3606 61436 3612
rect 60924 944 60976 950
rect 60924 886 60976 892
rect 62040 480 62068 3742
rect 63224 3256 63276 3262
rect 63224 3198 63276 3204
rect 63236 480 63264 3198
rect 63512 2106 63540 19774
rect 63788 15978 63816 19774
rect 63972 17610 64000 19774
rect 63960 17604 64012 17610
rect 63960 17546 64012 17552
rect 64156 16998 64184 19774
rect 64144 16992 64196 16998
rect 64144 16934 64196 16940
rect 64144 16652 64196 16658
rect 64144 16594 64196 16600
rect 63776 15972 63828 15978
rect 63776 15914 63828 15920
rect 63592 11824 63644 11830
rect 63592 11766 63644 11772
rect 63604 8265 63632 11766
rect 63590 8256 63646 8265
rect 63590 8191 63646 8200
rect 64156 3806 64184 16594
rect 64340 15094 64368 19774
rect 64524 16658 64552 19774
rect 64512 16652 64564 16658
rect 64512 16594 64564 16600
rect 64236 15088 64288 15094
rect 64236 15030 64288 15036
rect 64328 15088 64380 15094
rect 64328 15030 64380 15036
rect 64248 14618 64276 15030
rect 64236 14612 64288 14618
rect 64236 14554 64288 14560
rect 64708 14278 64736 19774
rect 64800 19774 64874 19802
rect 64984 19774 65058 19802
rect 65168 19774 65242 19802
rect 65352 19774 65426 19802
rect 65536 19774 65610 19802
rect 65766 19802 65794 20060
rect 65950 19802 65978 20060
rect 66134 19802 66162 20060
rect 65766 19774 65840 19802
rect 65950 19774 66024 19802
rect 64696 14272 64748 14278
rect 64696 14214 64748 14220
rect 64800 9994 64828 19774
rect 64984 18766 65012 19774
rect 64972 18760 65024 18766
rect 64972 18702 65024 18708
rect 65064 15700 65116 15706
rect 65064 15642 65116 15648
rect 64788 9988 64840 9994
rect 64788 9930 64840 9936
rect 64328 8900 64380 8906
rect 64328 8842 64380 8848
rect 64144 3800 64196 3806
rect 64144 3742 64196 3748
rect 63500 2100 63552 2106
rect 63500 2042 63552 2048
rect 64340 480 64368 8842
rect 64880 7744 64932 7750
rect 64880 7686 64932 7692
rect 64892 1222 64920 7686
rect 64880 1216 64932 1222
rect 64880 1158 64932 1164
rect 53300 354 53328 462
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 15642
rect 65168 14822 65196 19774
rect 65156 14816 65208 14822
rect 65156 14758 65208 14764
rect 65352 6118 65380 19774
rect 65536 18290 65564 19774
rect 65524 18284 65576 18290
rect 65524 18226 65576 18232
rect 65524 17536 65576 17542
rect 65524 17478 65576 17484
rect 65536 17134 65564 17478
rect 65524 17128 65576 17134
rect 65524 17070 65576 17076
rect 65708 17128 65760 17134
rect 65708 17070 65760 17076
rect 65616 16652 65668 16658
rect 65616 16594 65668 16600
rect 65524 15088 65576 15094
rect 65524 15030 65576 15036
rect 65536 11830 65564 15030
rect 65524 11824 65576 11830
rect 65524 11766 65576 11772
rect 65628 9246 65656 16594
rect 65720 13802 65748 17070
rect 65708 13796 65760 13802
rect 65708 13738 65760 13744
rect 65812 13462 65840 19774
rect 65892 17400 65944 17406
rect 65892 17342 65944 17348
rect 65904 17202 65932 17342
rect 65892 17196 65944 17202
rect 65892 17138 65944 17144
rect 65996 15366 66024 19774
rect 66088 19774 66162 19802
rect 66318 19802 66346 20060
rect 66502 19938 66530 20060
rect 66502 19910 66576 19938
rect 66444 19848 66496 19854
rect 66318 19774 66392 19802
rect 66444 19790 66496 19796
rect 66088 17746 66116 19774
rect 66076 17740 66128 17746
rect 66076 17682 66128 17688
rect 66076 17604 66128 17610
rect 66076 17546 66128 17552
rect 65984 15360 66036 15366
rect 65984 15302 66036 15308
rect 66088 15298 66116 17546
rect 66260 17400 66312 17406
rect 66260 17342 66312 17348
rect 66272 16522 66300 17342
rect 66364 16658 66392 19774
rect 66456 18494 66484 19790
rect 66444 18488 66496 18494
rect 66444 18430 66496 18436
rect 66444 16788 66496 16794
rect 66444 16730 66496 16736
rect 66352 16652 66404 16658
rect 66352 16594 66404 16600
rect 66260 16516 66312 16522
rect 66260 16458 66312 16464
rect 66168 15972 66220 15978
rect 66168 15914 66220 15920
rect 66260 15972 66312 15978
rect 66260 15914 66312 15920
rect 66076 15292 66128 15298
rect 66076 15234 66128 15240
rect 65800 13456 65852 13462
rect 65800 13398 65852 13404
rect 66180 10946 66208 15914
rect 66272 15774 66300 15914
rect 66260 15768 66312 15774
rect 66260 15710 66312 15716
rect 66456 13734 66484 16730
rect 66548 14074 66576 19910
rect 66686 19802 66714 20060
rect 66870 19802 66898 20060
rect 67054 19802 67082 20060
rect 67238 19802 67266 20060
rect 67422 19802 67450 20060
rect 67606 19802 67634 20060
rect 67790 19802 67818 20060
rect 67974 19802 68002 20060
rect 68158 19802 68186 20060
rect 68342 19802 68370 20060
rect 68526 19802 68554 20060
rect 66640 19774 66714 19802
rect 66824 19774 66898 19802
rect 67008 19774 67082 19802
rect 67192 19774 67266 19802
rect 67376 19774 67450 19802
rect 67560 19774 67634 19802
rect 67744 19774 67818 19802
rect 67928 19774 68002 19802
rect 68112 19774 68186 19802
rect 68296 19774 68370 19802
rect 68480 19774 68554 19802
rect 68710 19802 68738 20060
rect 68894 19802 68922 20060
rect 68710 19774 68784 19802
rect 66640 17814 66668 19774
rect 66628 17808 66680 17814
rect 66628 17750 66680 17756
rect 66824 16726 66852 19774
rect 66812 16720 66864 16726
rect 66812 16662 66864 16668
rect 66536 14068 66588 14074
rect 66536 14010 66588 14016
rect 66444 13728 66496 13734
rect 66444 13670 66496 13676
rect 66904 11960 66956 11966
rect 66904 11902 66956 11908
rect 66168 10940 66220 10946
rect 66168 10882 66220 10888
rect 65800 10600 65852 10606
rect 65800 10542 65852 10548
rect 65616 9240 65668 9246
rect 65616 9182 65668 9188
rect 65812 8226 65840 10542
rect 65800 8220 65852 8226
rect 65800 8162 65852 8168
rect 65340 6112 65392 6118
rect 65340 6054 65392 6060
rect 66720 5160 66772 5166
rect 66720 5102 66772 5108
rect 66732 480 66760 5102
rect 66916 3602 66944 11902
rect 67008 5846 67036 19774
rect 67192 18834 67220 19774
rect 67180 18828 67232 18834
rect 67180 18770 67232 18776
rect 67376 12306 67404 19774
rect 67364 12300 67416 12306
rect 67364 12242 67416 12248
rect 67560 11422 67588 19774
rect 67744 17882 67772 19774
rect 67732 17876 67784 17882
rect 67732 17818 67784 17824
rect 67732 17740 67784 17746
rect 67732 17682 67784 17688
rect 67638 15872 67694 15881
rect 67638 15807 67694 15816
rect 67652 13802 67680 15807
rect 67744 14618 67772 17682
rect 67824 16856 67876 16862
rect 67824 16798 67876 16804
rect 67732 14612 67784 14618
rect 67732 14554 67784 14560
rect 67640 13796 67692 13802
rect 67640 13738 67692 13744
rect 67836 13666 67864 16798
rect 67928 16794 67956 19774
rect 67916 16788 67968 16794
rect 67916 16730 67968 16736
rect 67824 13660 67876 13666
rect 67824 13602 67876 13608
rect 67640 11892 67692 11898
rect 67640 11834 67692 11840
rect 67548 11416 67600 11422
rect 67548 11358 67600 11364
rect 66996 5840 67048 5846
rect 66996 5782 67048 5788
rect 67548 5568 67600 5574
rect 67548 5510 67600 5516
rect 66904 3596 66956 3602
rect 66904 3538 66956 3544
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67560 66 67588 5510
rect 67652 354 67680 11834
rect 67916 9104 67968 9110
rect 67916 9046 67968 9052
rect 67928 2378 67956 9046
rect 68112 8566 68140 19774
rect 68296 17678 68324 19774
rect 68284 17672 68336 17678
rect 68284 17614 68336 17620
rect 68376 17672 68428 17678
rect 68376 17614 68428 17620
rect 68284 16652 68336 16658
rect 68284 16594 68336 16600
rect 68296 8634 68324 16594
rect 68388 13598 68416 17614
rect 68376 13592 68428 13598
rect 68376 13534 68428 13540
rect 68480 10878 68508 19774
rect 68756 13054 68784 19774
rect 68848 19774 68922 19802
rect 69078 19802 69106 20060
rect 69262 19802 69290 20060
rect 69446 19802 69474 20060
rect 69630 19802 69658 20060
rect 69078 19774 69152 19802
rect 69262 19774 69336 19802
rect 68848 18358 68876 19774
rect 68836 18352 68888 18358
rect 68836 18294 68888 18300
rect 68836 13116 68888 13122
rect 68836 13058 68888 13064
rect 68744 13048 68796 13054
rect 68744 12990 68796 12996
rect 68468 10872 68520 10878
rect 68468 10814 68520 10820
rect 68560 10464 68612 10470
rect 68560 10406 68612 10412
rect 68284 8628 68336 8634
rect 68284 8570 68336 8576
rect 68100 8560 68152 8566
rect 68100 8502 68152 8508
rect 68572 4826 68600 10406
rect 68652 10396 68704 10402
rect 68652 10338 68704 10344
rect 68560 4820 68612 4826
rect 68560 4762 68612 4768
rect 68664 4690 68692 10338
rect 68744 9988 68796 9994
rect 68744 9930 68796 9936
rect 68756 6186 68784 9930
rect 68848 9110 68876 13058
rect 68928 10396 68980 10402
rect 68928 10338 68980 10344
rect 68940 9586 68968 10338
rect 68928 9580 68980 9586
rect 68928 9522 68980 9528
rect 68836 9104 68888 9110
rect 68836 9046 68888 9052
rect 69124 7070 69152 19774
rect 69308 17610 69336 19774
rect 69400 19774 69474 19802
rect 69584 19774 69658 19802
rect 69814 19802 69842 20060
rect 69998 19802 70026 20060
rect 70182 19802 70210 20060
rect 70366 19802 70394 20060
rect 70550 19802 70578 20060
rect 70734 19802 70762 20060
rect 70918 19802 70946 20060
rect 71102 19802 71130 20060
rect 71286 19802 71314 20060
rect 71470 19802 71498 20060
rect 71654 19802 71682 20060
rect 69814 19774 69888 19802
rect 69400 19174 69428 19774
rect 69388 19168 69440 19174
rect 69388 19110 69440 19116
rect 69296 17604 69348 17610
rect 69296 17546 69348 17552
rect 69584 12374 69612 19774
rect 69860 14754 69888 19774
rect 69952 19774 70026 19802
rect 70136 19774 70210 19802
rect 70320 19774 70394 19802
rect 70504 19774 70578 19802
rect 70688 19774 70762 19802
rect 70872 19774 70946 19802
rect 71056 19774 71130 19802
rect 71240 19774 71314 19802
rect 71424 19774 71498 19802
rect 71608 19774 71682 19802
rect 71838 19802 71866 20060
rect 72022 19802 72050 20060
rect 72206 19802 72234 20060
rect 72390 19802 72418 20060
rect 71838 19774 71912 19802
rect 69952 18562 69980 19774
rect 69940 18556 69992 18562
rect 69940 18498 69992 18504
rect 70136 16862 70164 19774
rect 70124 16856 70176 16862
rect 70124 16798 70176 16804
rect 69848 14748 69900 14754
rect 69848 14690 69900 14696
rect 69848 14204 69900 14210
rect 69848 14146 69900 14152
rect 69572 12368 69624 12374
rect 69572 12310 69624 12316
rect 69112 7064 69164 7070
rect 69112 7006 69164 7012
rect 69112 6588 69164 6594
rect 69112 6530 69164 6536
rect 68744 6180 68796 6186
rect 68744 6122 68796 6128
rect 68652 4684 68704 4690
rect 68652 4626 68704 4632
rect 67916 2372 67968 2378
rect 67916 2314 67968 2320
rect 69124 480 69152 6530
rect 69664 3800 69716 3806
rect 69664 3742 69716 3748
rect 69676 1018 69704 3742
rect 69664 1012 69716 1018
rect 69664 954 69716 960
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67548 60 67600 66
rect 67548 2 67600 8
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 14146
rect 70320 12306 70348 19774
rect 70504 16590 70532 19774
rect 70688 19718 70716 19774
rect 70676 19712 70728 19718
rect 70676 19654 70728 19660
rect 70584 18352 70636 18358
rect 70584 18294 70636 18300
rect 70492 16584 70544 16590
rect 70492 16526 70544 16532
rect 70492 15292 70544 15298
rect 70492 15234 70544 15240
rect 70400 13456 70452 13462
rect 70400 13398 70452 13404
rect 70308 12300 70360 12306
rect 70308 12242 70360 12248
rect 70412 9994 70440 13398
rect 70400 9988 70452 9994
rect 70400 9930 70452 9936
rect 70504 8906 70532 15234
rect 70596 11014 70624 18294
rect 70674 15872 70730 15881
rect 70674 15807 70730 15816
rect 70584 11008 70636 11014
rect 70584 10950 70636 10956
rect 70688 9518 70716 15807
rect 70872 12714 70900 19774
rect 71056 16318 71084 19774
rect 71240 18358 71268 19774
rect 71228 18352 71280 18358
rect 71228 18294 71280 18300
rect 71044 16312 71096 16318
rect 71044 16254 71096 16260
rect 71424 14890 71452 19774
rect 71608 17406 71636 19774
rect 71596 17400 71648 17406
rect 71596 17342 71648 17348
rect 71884 17066 71912 19774
rect 71976 19774 72050 19802
rect 72160 19774 72234 19802
rect 72344 19774 72418 19802
rect 72574 19802 72602 20060
rect 72758 19802 72786 20060
rect 72942 19802 72970 20060
rect 73126 19802 73154 20060
rect 72574 19774 72648 19802
rect 71872 17060 71924 17066
rect 71872 17002 71924 17008
rect 71780 16720 71832 16726
rect 71780 16662 71832 16668
rect 71792 15201 71820 16662
rect 71872 16312 71924 16318
rect 71872 16254 71924 16260
rect 71778 15192 71834 15201
rect 71778 15127 71834 15136
rect 71412 14884 71464 14890
rect 71412 14826 71464 14832
rect 71780 13796 71832 13802
rect 71780 13738 71832 13744
rect 70952 13388 71004 13394
rect 70952 13330 71004 13336
rect 70860 12708 70912 12714
rect 70860 12650 70912 12656
rect 70676 9512 70728 9518
rect 70676 9454 70728 9460
rect 70492 8900 70544 8906
rect 70492 8842 70544 8848
rect 70676 7948 70728 7954
rect 70676 7890 70728 7896
rect 70688 6089 70716 7890
rect 70674 6080 70730 6089
rect 70674 6015 70730 6024
rect 70964 3482 70992 13330
rect 71792 11490 71820 13738
rect 71688 11484 71740 11490
rect 71688 11426 71740 11432
rect 71780 11484 71832 11490
rect 71780 11426 71832 11432
rect 71700 11370 71728 11426
rect 71884 11370 71912 16254
rect 71700 11342 71912 11370
rect 71136 10940 71188 10946
rect 71136 10882 71188 10888
rect 71044 8220 71096 8226
rect 71044 8162 71096 8168
rect 71056 4865 71084 8162
rect 71042 4856 71098 4865
rect 71042 4791 71098 4800
rect 71148 3942 71176 10882
rect 71780 9036 71832 9042
rect 71780 8978 71832 8984
rect 71792 8129 71820 8978
rect 71778 8120 71834 8129
rect 71778 8055 71834 8064
rect 71976 5370 72004 19774
rect 72160 17202 72188 19774
rect 72148 17196 72200 17202
rect 72148 17138 72200 17144
rect 71964 5364 72016 5370
rect 71964 5306 72016 5312
rect 71136 3936 71188 3942
rect 71136 3878 71188 3884
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72344 1086 72372 19774
rect 72424 16652 72476 16658
rect 72424 16594 72476 16600
rect 72436 9654 72464 16594
rect 72620 12238 72648 19774
rect 72712 19774 72786 19802
rect 72896 19774 72970 19802
rect 73080 19774 73154 19802
rect 73310 19802 73338 20060
rect 73494 19802 73522 20060
rect 73678 19802 73706 20060
rect 73862 19802 73890 20060
rect 74046 19802 74074 20060
rect 74230 19802 74258 20060
rect 74414 19802 74442 20060
rect 74598 19802 74626 20060
rect 74782 19802 74810 20060
rect 73310 19774 73384 19802
rect 73494 19774 73568 19802
rect 72712 16930 72740 19774
rect 72700 16924 72752 16930
rect 72700 16866 72752 16872
rect 72608 12232 72660 12238
rect 72608 12174 72660 12180
rect 72424 9648 72476 9654
rect 72424 9590 72476 9596
rect 72896 6798 72924 19774
rect 73080 13666 73108 19774
rect 73356 16930 73384 19774
rect 73540 18834 73568 19774
rect 73632 19774 73706 19802
rect 73816 19774 73890 19802
rect 74000 19774 74074 19802
rect 74184 19774 74258 19802
rect 74368 19774 74442 19802
rect 74552 19774 74626 19802
rect 74736 19774 74810 19802
rect 74966 19802 74994 20060
rect 75150 19802 75178 20060
rect 75334 19802 75362 20060
rect 75518 19802 75546 20060
rect 75702 19802 75730 20060
rect 75886 19802 75914 20060
rect 76070 19802 76098 20060
rect 76254 19802 76282 20060
rect 76438 19802 76466 20060
rect 76622 19802 76650 20060
rect 76806 19802 76834 20060
rect 74966 19774 75040 19802
rect 73528 18828 73580 18834
rect 73528 18770 73580 18776
rect 73344 16924 73396 16930
rect 73344 16866 73396 16872
rect 73632 15774 73660 19774
rect 73816 18698 73844 19774
rect 73804 18692 73856 18698
rect 73804 18634 73856 18640
rect 73896 17468 73948 17474
rect 73896 17410 73948 17416
rect 73804 16244 73856 16250
rect 73804 16186 73856 16192
rect 73620 15768 73672 15774
rect 73620 15710 73672 15716
rect 73068 13660 73120 13666
rect 73068 13602 73120 13608
rect 72884 6792 72936 6798
rect 72884 6734 72936 6740
rect 72608 6520 72660 6526
rect 72608 6462 72660 6468
rect 72332 1080 72384 1086
rect 72332 1022 72384 1028
rect 72620 480 72648 6462
rect 73816 5386 73844 16186
rect 73908 6526 73936 17410
rect 74000 17134 74028 19774
rect 73988 17128 74040 17134
rect 73988 17070 74040 17076
rect 73896 6520 73948 6526
rect 73896 6462 73948 6468
rect 73816 5358 73936 5386
rect 73804 4752 73856 4758
rect 73804 4694 73856 4700
rect 73816 480 73844 4694
rect 73908 3806 73936 5358
rect 74184 5234 74212 19774
rect 74172 5228 74224 5234
rect 74172 5170 74224 5176
rect 73896 3800 73948 3806
rect 73896 3742 73948 3748
rect 74368 2038 74396 19774
rect 74552 16182 74580 19774
rect 74540 16176 74592 16182
rect 74540 16118 74592 16124
rect 74736 7954 74764 19774
rect 75012 19174 75040 19774
rect 75104 19774 75178 19802
rect 75288 19774 75362 19802
rect 75472 19774 75546 19802
rect 75656 19774 75730 19802
rect 75840 19774 75914 19802
rect 76024 19774 76098 19802
rect 76208 19774 76282 19802
rect 76392 19774 76466 19802
rect 76576 19774 76650 19802
rect 76760 19774 76834 19802
rect 76990 19802 77018 20060
rect 77174 19802 77202 20060
rect 77358 19802 77386 20060
rect 77542 19802 77570 20060
rect 76990 19774 77064 19802
rect 75000 19168 75052 19174
rect 75000 19110 75052 19116
rect 75104 17406 75132 19774
rect 75184 17536 75236 17542
rect 75184 17478 75236 17484
rect 75092 17400 75144 17406
rect 75092 17342 75144 17348
rect 75000 13320 75052 13326
rect 75000 13262 75052 13268
rect 74724 7948 74776 7954
rect 74724 7890 74776 7896
rect 74356 2032 74408 2038
rect 74356 1974 74408 1980
rect 75012 480 75040 13262
rect 75196 4146 75224 17478
rect 75288 13734 75316 19774
rect 75276 13728 75328 13734
rect 75276 13670 75328 13676
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 75472 1970 75500 19774
rect 75656 15230 75684 19774
rect 75644 15224 75696 15230
rect 75644 15166 75696 15172
rect 75840 12170 75868 19774
rect 75828 12164 75880 12170
rect 75828 12106 75880 12112
rect 75920 10736 75972 10742
rect 75920 10678 75972 10684
rect 75460 1964 75512 1970
rect 75460 1906 75512 1912
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 10678
rect 76024 2446 76052 19774
rect 76104 18624 76156 18630
rect 76104 18566 76156 18572
rect 76116 14793 76144 18566
rect 76102 14784 76158 14793
rect 76102 14719 76158 14728
rect 76208 4622 76236 19774
rect 76392 14686 76420 19774
rect 76380 14680 76432 14686
rect 76380 14622 76432 14628
rect 76196 4616 76248 4622
rect 76196 4558 76248 4564
rect 76576 2718 76604 19774
rect 76760 16658 76788 19774
rect 77036 17678 77064 19774
rect 77128 19774 77202 19802
rect 77312 19774 77386 19802
rect 77496 19774 77570 19802
rect 77726 19802 77754 20060
rect 77910 19802 77938 20060
rect 77726 19774 77800 19802
rect 77024 17672 77076 17678
rect 77024 17614 77076 17620
rect 76748 16652 76800 16658
rect 76748 16594 76800 16600
rect 77024 16176 77076 16182
rect 77024 16118 77076 16124
rect 77036 11354 77064 16118
rect 77024 11348 77076 11354
rect 77024 11290 77076 11296
rect 76564 2712 76616 2718
rect 76564 2654 76616 2660
rect 76012 2440 76064 2446
rect 76012 2382 76064 2388
rect 77128 1154 77156 19774
rect 77312 15162 77340 19774
rect 77300 15156 77352 15162
rect 77300 15098 77352 15104
rect 77208 14136 77260 14142
rect 77208 14078 77260 14084
rect 77220 11966 77248 14078
rect 77496 13122 77524 19774
rect 77772 18630 77800 19774
rect 77864 19774 77938 19802
rect 78094 19802 78122 20060
rect 78278 19802 78306 20060
rect 78462 19802 78490 20060
rect 78646 19802 78674 20060
rect 78830 19802 78858 20060
rect 79014 19802 79042 20060
rect 79198 19802 79226 20060
rect 79382 19802 79410 20060
rect 79566 19802 79594 20060
rect 79750 19802 79778 20060
rect 78094 19774 78168 19802
rect 77760 18624 77812 18630
rect 77760 18566 77812 18572
rect 77864 15434 77892 19774
rect 78140 17202 78168 19774
rect 78232 19774 78306 19802
rect 78416 19774 78490 19802
rect 78600 19774 78674 19802
rect 78784 19774 78858 19802
rect 78968 19774 79042 19802
rect 79152 19774 79226 19802
rect 79336 19774 79410 19802
rect 79520 19774 79594 19802
rect 79704 19774 79778 19802
rect 79934 19802 79962 20060
rect 80118 19802 80146 20060
rect 79934 19774 80008 19802
rect 78128 17196 78180 17202
rect 78128 17138 78180 17144
rect 77852 15428 77904 15434
rect 77852 15370 77904 15376
rect 77484 13116 77536 13122
rect 77484 13058 77536 13064
rect 77208 11960 77260 11966
rect 77208 11902 77260 11908
rect 77208 11756 77260 11762
rect 77208 11698 77260 11704
rect 77220 10849 77248 11698
rect 77206 10840 77262 10849
rect 77206 10775 77262 10784
rect 78128 10192 78180 10198
rect 78128 10134 78180 10140
rect 77392 5024 77444 5030
rect 77392 4966 77444 4972
rect 77116 1148 77168 1154
rect 77116 1090 77168 1096
rect 77404 480 77432 4966
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10134
rect 78232 2582 78260 19774
rect 78312 14748 78364 14754
rect 78312 14690 78364 14696
rect 78324 8362 78352 14690
rect 78416 10946 78444 19774
rect 78496 15224 78548 15230
rect 78496 15166 78548 15172
rect 78508 13598 78536 15166
rect 78496 13592 78548 13598
rect 78496 13534 78548 13540
rect 78404 10940 78456 10946
rect 78404 10882 78456 10888
rect 78600 10198 78628 19774
rect 78680 13864 78732 13870
rect 78680 13806 78732 13812
rect 78692 12102 78720 13806
rect 78680 12096 78732 12102
rect 78680 12038 78732 12044
rect 78588 10192 78640 10198
rect 78588 10134 78640 10140
rect 78312 8356 78364 8362
rect 78312 8298 78364 8304
rect 78220 2576 78272 2582
rect 78220 2518 78272 2524
rect 78784 610 78812 19774
rect 78968 14006 78996 19774
rect 79152 17610 79180 19774
rect 79140 17604 79192 17610
rect 79140 17546 79192 17552
rect 79140 14612 79192 14618
rect 79140 14554 79192 14560
rect 78956 14000 79008 14006
rect 78956 13942 79008 13948
rect 79152 11762 79180 14554
rect 79232 14544 79284 14550
rect 79232 14486 79284 14492
rect 79244 14210 79272 14486
rect 79232 14204 79284 14210
rect 79232 14146 79284 14152
rect 79232 13184 79284 13190
rect 79232 13126 79284 13132
rect 79140 11756 79192 11762
rect 79140 11698 79192 11704
rect 79244 10713 79272 13126
rect 79230 10704 79286 10713
rect 79230 10639 79286 10648
rect 78772 604 78824 610
rect 78772 546 78824 552
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79336 134 79364 19774
rect 79416 17672 79468 17678
rect 79416 17614 79468 17620
rect 79428 5302 79456 17614
rect 79520 16318 79548 19774
rect 79508 16312 79560 16318
rect 79508 16254 79560 16260
rect 79508 14476 79560 14482
rect 79508 14418 79560 14424
rect 79416 5296 79468 5302
rect 79416 5238 79468 5244
rect 79520 3398 79548 14418
rect 79704 14142 79732 19774
rect 79980 18358 80008 19774
rect 80072 19774 80146 19802
rect 80302 19802 80330 20060
rect 80486 19802 80514 20060
rect 80670 19802 80698 20060
rect 80854 19802 80882 20060
rect 80302 19774 80376 19802
rect 80486 19774 80560 19802
rect 79968 18352 80020 18358
rect 79968 18294 80020 18300
rect 79692 14136 79744 14142
rect 79692 14078 79744 14084
rect 79692 6452 79744 6458
rect 79692 6394 79744 6400
rect 79508 3392 79560 3398
rect 79508 3334 79560 3340
rect 79704 480 79732 6394
rect 80072 5982 80100 19774
rect 80150 18728 80206 18737
rect 80150 18663 80206 18672
rect 80164 17377 80192 18663
rect 80348 17950 80376 19774
rect 80532 18766 80560 19774
rect 80624 19774 80698 19802
rect 80808 19774 80882 19802
rect 81038 19802 81066 20060
rect 81222 19802 81250 20060
rect 81406 19802 81434 20060
rect 81590 19802 81618 20060
rect 81774 19802 81802 20060
rect 81958 19802 81986 20060
rect 81038 19774 81112 19802
rect 80520 18760 80572 18766
rect 80520 18702 80572 18708
rect 80336 17944 80388 17950
rect 80336 17886 80388 17892
rect 80150 17368 80206 17377
rect 80150 17303 80206 17312
rect 80624 8158 80652 19774
rect 80704 17400 80756 17406
rect 80704 17342 80756 17348
rect 80612 8152 80664 8158
rect 80612 8094 80664 8100
rect 80612 6180 80664 6186
rect 80612 6122 80664 6128
rect 80060 5976 80112 5982
rect 80060 5918 80112 5924
rect 80624 3777 80652 6122
rect 80610 3768 80666 3777
rect 80610 3703 80666 3712
rect 80716 1834 80744 17342
rect 80808 13394 80836 19774
rect 81084 17406 81112 19774
rect 81176 19774 81250 19802
rect 81360 19774 81434 19802
rect 81544 19774 81618 19802
rect 81728 19774 81802 19802
rect 81912 19774 81986 19802
rect 82142 19802 82170 20060
rect 82326 19802 82354 20060
rect 82510 19802 82538 20060
rect 82142 19774 82216 19802
rect 81072 17400 81124 17406
rect 81072 17342 81124 17348
rect 80888 14000 80940 14006
rect 80888 13942 80940 13948
rect 80796 13388 80848 13394
rect 80796 13330 80848 13336
rect 80900 9518 80928 13942
rect 81176 13530 81204 19774
rect 81360 15230 81388 19774
rect 81440 19712 81492 19718
rect 81440 19654 81492 19660
rect 81452 19310 81480 19654
rect 81440 19304 81492 19310
rect 81440 19246 81492 19252
rect 81440 17944 81492 17950
rect 81440 17886 81492 17892
rect 81452 15858 81480 17886
rect 81544 16182 81572 19774
rect 81624 16788 81676 16794
rect 81624 16730 81676 16736
rect 81532 16176 81584 16182
rect 81532 16118 81584 16124
rect 81452 15830 81572 15858
rect 81440 15768 81492 15774
rect 81440 15710 81492 15716
rect 81348 15224 81400 15230
rect 81348 15166 81400 15172
rect 81452 14822 81480 15710
rect 81440 14816 81492 14822
rect 81440 14758 81492 14764
rect 81544 14482 81572 15830
rect 81532 14476 81584 14482
rect 81532 14418 81584 14424
rect 81440 14068 81492 14074
rect 81440 14010 81492 14016
rect 81164 13524 81216 13530
rect 81164 13466 81216 13472
rect 81452 12374 81480 14010
rect 81440 12368 81492 12374
rect 81440 12310 81492 12316
rect 81532 11960 81584 11966
rect 81532 11902 81584 11908
rect 81348 11824 81400 11830
rect 81348 11766 81400 11772
rect 80888 9512 80940 9518
rect 80888 9454 80940 9460
rect 81360 8226 81388 11766
rect 81544 9042 81572 11902
rect 81636 9926 81664 16730
rect 81728 15502 81756 19774
rect 81716 15496 81768 15502
rect 81716 15438 81768 15444
rect 81912 14754 81940 19774
rect 82188 18698 82216 19774
rect 82280 19774 82354 19802
rect 82464 19774 82538 19802
rect 82694 19802 82722 20060
rect 82878 19802 82906 20060
rect 83062 19802 83090 20060
rect 83246 19802 83274 20060
rect 83430 19802 83458 20060
rect 83614 19802 83642 20060
rect 82694 19774 82768 19802
rect 82878 19774 82952 19802
rect 82176 18692 82228 18698
rect 82176 18634 82228 18640
rect 81992 17536 82044 17542
rect 81992 17478 82044 17484
rect 81900 14748 81952 14754
rect 81900 14690 81952 14696
rect 82004 13870 82032 17478
rect 82176 17468 82228 17474
rect 82176 17410 82228 17416
rect 82188 14006 82216 17410
rect 82176 14000 82228 14006
rect 82176 13942 82228 13948
rect 81992 13864 82044 13870
rect 81992 13806 82044 13812
rect 82176 13252 82228 13258
rect 82176 13194 82228 13200
rect 81624 9920 81676 9926
rect 81624 9862 81676 9868
rect 81532 9036 81584 9042
rect 81532 8978 81584 8984
rect 82084 8968 82136 8974
rect 82084 8910 82136 8916
rect 81348 8220 81400 8226
rect 81348 8162 81400 8168
rect 81348 7676 81400 7682
rect 81348 7618 81400 7624
rect 80888 7608 80940 7614
rect 80888 7550 80940 7556
rect 80900 6730 80928 7550
rect 80888 6724 80940 6730
rect 80888 6666 80940 6672
rect 81360 5137 81388 7618
rect 82096 6633 82124 8910
rect 82082 6624 82138 6633
rect 82082 6559 82138 6568
rect 82084 6520 82136 6526
rect 82084 6462 82136 6468
rect 81346 5128 81402 5137
rect 80888 5092 80940 5098
rect 81346 5063 81402 5072
rect 80888 5034 80940 5040
rect 80704 1828 80756 1834
rect 80704 1770 80756 1776
rect 80900 480 80928 5034
rect 81440 3528 81492 3534
rect 81440 3470 81492 3476
rect 81452 2242 81480 3470
rect 81440 2236 81492 2242
rect 81440 2178 81492 2184
rect 82096 480 82124 6462
rect 82188 3262 82216 13194
rect 82280 10742 82308 19774
rect 82360 17196 82412 17202
rect 82360 17138 82412 17144
rect 82372 11966 82400 17138
rect 82464 16182 82492 19774
rect 82740 17882 82768 19774
rect 82820 19644 82872 19650
rect 82820 19586 82872 19592
rect 82728 17876 82780 17882
rect 82728 17818 82780 17824
rect 82832 16998 82860 19586
rect 82820 16992 82872 16998
rect 82820 16934 82872 16940
rect 82924 16726 82952 19774
rect 83016 19774 83090 19802
rect 83200 19774 83274 19802
rect 83384 19774 83458 19802
rect 83568 19774 83642 19802
rect 83798 19802 83826 20060
rect 83982 19802 84010 20060
rect 84166 19802 84194 20060
rect 84350 19802 84378 20060
rect 84534 19802 84562 20060
rect 84718 19802 84746 20060
rect 83798 19774 83872 19802
rect 82912 16720 82964 16726
rect 82912 16662 82964 16668
rect 82452 16176 82504 16182
rect 82452 16118 82504 16124
rect 82544 15224 82596 15230
rect 82544 15166 82596 15172
rect 82360 11960 82412 11966
rect 82360 11902 82412 11908
rect 82556 11898 82584 15166
rect 82544 11892 82596 11898
rect 82544 11834 82596 11840
rect 82450 11792 82506 11801
rect 82450 11727 82506 11736
rect 82268 10736 82320 10742
rect 82268 10678 82320 10684
rect 82464 10402 82492 11727
rect 82728 11552 82780 11558
rect 82728 11494 82780 11500
rect 82452 10396 82504 10402
rect 82452 10338 82504 10344
rect 82740 8770 82768 11494
rect 82728 8764 82780 8770
rect 82728 8706 82780 8712
rect 83016 5166 83044 19774
rect 83200 13802 83228 19774
rect 83188 13796 83240 13802
rect 83188 13738 83240 13744
rect 83186 11656 83242 11665
rect 83186 11591 83242 11600
rect 83200 5506 83228 11591
rect 83280 9376 83332 9382
rect 83280 9318 83332 9324
rect 83188 5500 83240 5506
rect 83188 5442 83240 5448
rect 83004 5160 83056 5166
rect 83004 5102 83056 5108
rect 82176 3256 82228 3262
rect 82176 3198 82228 3204
rect 83292 480 83320 9318
rect 83384 8838 83412 19774
rect 83568 10402 83596 19774
rect 83844 16998 83872 19774
rect 83936 19774 84010 19802
rect 84120 19774 84194 19802
rect 84304 19774 84378 19802
rect 84488 19774 84562 19802
rect 84672 19774 84746 19802
rect 84902 19802 84930 20060
rect 85086 19802 85114 20060
rect 85270 19802 85298 20060
rect 85454 19802 85482 20060
rect 85638 19802 85666 20060
rect 84902 19774 84976 19802
rect 83832 16992 83884 16998
rect 83832 16934 83884 16940
rect 83936 16522 83964 19774
rect 83924 16516 83976 16522
rect 83924 16458 83976 16464
rect 84120 15638 84148 19774
rect 84304 17474 84332 19774
rect 84384 19032 84436 19038
rect 84384 18974 84436 18980
rect 84292 17468 84344 17474
rect 84292 17410 84344 17416
rect 84108 15632 84160 15638
rect 84108 15574 84160 15580
rect 84396 11937 84424 18974
rect 84488 16794 84516 19774
rect 84476 16788 84528 16794
rect 84476 16730 84528 16736
rect 84672 12850 84700 19774
rect 84948 18426 84976 19774
rect 85040 19774 85114 19802
rect 85224 19774 85298 19802
rect 85408 19774 85482 19802
rect 85592 19774 85666 19802
rect 85822 19802 85850 20060
rect 86006 19802 86034 20060
rect 86190 19802 86218 20060
rect 86374 19802 86402 20060
rect 85822 19774 85896 19802
rect 84936 18420 84988 18426
rect 84936 18362 84988 18368
rect 84844 16992 84896 16998
rect 84844 16934 84896 16940
rect 84660 12844 84712 12850
rect 84660 12786 84712 12792
rect 84382 11928 84438 11937
rect 84382 11863 84438 11872
rect 84568 11484 84620 11490
rect 84568 11426 84620 11432
rect 83556 10396 83608 10402
rect 83556 10338 83608 10344
rect 84580 9722 84608 11426
rect 84568 9716 84620 9722
rect 84568 9658 84620 9664
rect 84752 9240 84804 9246
rect 84752 9182 84804 9188
rect 83372 8832 83424 8838
rect 83372 8774 83424 8780
rect 84660 8832 84712 8838
rect 84660 8774 84712 8780
rect 84384 8356 84436 8362
rect 84384 8298 84436 8304
rect 84396 5438 84424 8298
rect 84384 5432 84436 5438
rect 84384 5374 84436 5380
rect 84672 5098 84700 8774
rect 84764 7410 84792 9182
rect 84752 7404 84804 7410
rect 84752 7346 84804 7352
rect 84660 5092 84712 5098
rect 84660 5034 84712 5040
rect 84476 4956 84528 4962
rect 84476 4898 84528 4904
rect 84488 480 84516 4898
rect 84856 746 84884 16934
rect 84936 14204 84988 14210
rect 84936 14146 84988 14152
rect 84948 3330 84976 14146
rect 85040 12102 85068 19774
rect 85120 16720 85172 16726
rect 85120 16662 85172 16668
rect 85028 12096 85080 12102
rect 85028 12038 85080 12044
rect 85028 8220 85080 8226
rect 85028 8162 85080 8168
rect 85040 4010 85068 8162
rect 85132 6662 85160 16662
rect 85224 8974 85252 19774
rect 85408 18494 85436 19774
rect 85396 18488 85448 18494
rect 85396 18430 85448 18436
rect 85488 18148 85540 18154
rect 85488 18090 85540 18096
rect 85500 16930 85528 18090
rect 85488 16924 85540 16930
rect 85488 16866 85540 16872
rect 85212 8968 85264 8974
rect 85212 8910 85264 8916
rect 85120 6656 85172 6662
rect 85120 6598 85172 6604
rect 85592 6594 85620 19774
rect 85764 18080 85816 18086
rect 85764 18022 85816 18028
rect 85776 10810 85804 18022
rect 85868 16862 85896 19774
rect 85960 19774 86034 19802
rect 86144 19774 86218 19802
rect 86328 19774 86402 19802
rect 86558 19802 86586 20060
rect 86742 19802 86770 20060
rect 86926 19802 86954 20060
rect 86558 19774 86632 19802
rect 85856 16856 85908 16862
rect 85856 16798 85908 16804
rect 85764 10804 85816 10810
rect 85764 10746 85816 10752
rect 85580 6588 85632 6594
rect 85580 6530 85632 6536
rect 85028 4004 85080 4010
rect 85028 3946 85080 3952
rect 85672 3868 85724 3874
rect 85672 3810 85724 3816
rect 84936 3324 84988 3330
rect 84936 3266 84988 3272
rect 84844 740 84896 746
rect 84844 682 84896 688
rect 85684 480 85712 3810
rect 85960 1290 85988 19774
rect 86144 14618 86172 19774
rect 86132 14612 86184 14618
rect 86132 14554 86184 14560
rect 86328 6458 86356 19774
rect 86604 17678 86632 19774
rect 86696 19774 86770 19802
rect 86880 19774 86954 19802
rect 87110 19802 87138 20060
rect 87294 19802 87322 20060
rect 87110 19774 87184 19802
rect 86592 17672 86644 17678
rect 86592 17614 86644 17620
rect 86500 16516 86552 16522
rect 86500 16458 86552 16464
rect 86512 9382 86540 16458
rect 86696 13326 86724 19774
rect 86776 18964 86828 18970
rect 86776 18906 86828 18912
rect 86788 17950 86816 18906
rect 86776 17944 86828 17950
rect 86776 17886 86828 17892
rect 86776 13796 86828 13802
rect 86776 13738 86828 13744
rect 86684 13320 86736 13326
rect 86684 13262 86736 13268
rect 86788 9654 86816 13738
rect 86776 9648 86828 9654
rect 86776 9590 86828 9596
rect 86500 9376 86552 9382
rect 86500 9318 86552 9324
rect 86880 8650 86908 19774
rect 87156 18737 87184 19774
rect 87248 19774 87322 19802
rect 87478 19802 87506 20060
rect 87662 19802 87690 20060
rect 87846 19802 87874 20060
rect 87478 19774 87552 19802
rect 87662 19774 87736 19802
rect 87142 18728 87198 18737
rect 87142 18663 87198 18672
rect 86960 16108 87012 16114
rect 86960 16050 87012 16056
rect 86972 15298 87000 16050
rect 86960 15292 87012 15298
rect 86960 15234 87012 15240
rect 86960 9104 87012 9110
rect 86960 9046 87012 9052
rect 86788 8622 86908 8650
rect 86316 6452 86368 6458
rect 86316 6394 86368 6400
rect 86684 5500 86736 5506
rect 86684 5442 86736 5448
rect 86696 2553 86724 5442
rect 86788 4962 86816 8622
rect 86972 7993 87000 9046
rect 86958 7984 87014 7993
rect 86958 7919 87014 7928
rect 87248 6526 87276 19774
rect 87524 17610 87552 19774
rect 87708 18970 87736 19774
rect 87800 19774 87874 19802
rect 88030 19802 88058 20060
rect 88214 19802 88242 20060
rect 88398 19802 88426 20060
rect 88582 19802 88610 20060
rect 88766 19802 88794 20060
rect 88950 19802 88978 20060
rect 89134 19802 89162 20060
rect 89318 19802 89346 20060
rect 89502 19802 89530 20060
rect 89686 19802 89714 20060
rect 89870 19802 89898 20060
rect 90054 19802 90082 20060
rect 90238 19802 90266 20060
rect 90422 19802 90450 20060
rect 90606 19802 90634 20060
rect 88030 19774 88104 19802
rect 88214 19774 88288 19802
rect 87696 18964 87748 18970
rect 87696 18906 87748 18912
rect 87512 17604 87564 17610
rect 87512 17546 87564 17552
rect 87604 17400 87656 17406
rect 87604 17342 87656 17348
rect 87236 6520 87288 6526
rect 87236 6462 87288 6468
rect 86868 6384 86920 6390
rect 86868 6326 86920 6332
rect 86776 4956 86828 4962
rect 86776 4898 86828 4904
rect 86682 2544 86738 2553
rect 86682 2479 86738 2488
rect 85948 1284 86000 1290
rect 85948 1226 86000 1232
rect 86880 480 86908 6326
rect 86960 6248 87012 6254
rect 86960 6190 87012 6196
rect 86972 5506 87000 6190
rect 86960 5500 87012 5506
rect 86960 5442 87012 5448
rect 87616 2310 87644 17342
rect 87696 16176 87748 16182
rect 87696 16118 87748 16124
rect 87708 6186 87736 16118
rect 87800 15230 87828 19774
rect 87972 19440 88024 19446
rect 87972 19382 88024 19388
rect 87984 18086 88012 19382
rect 87972 18080 88024 18086
rect 87972 18022 88024 18028
rect 88076 17746 88104 19774
rect 88064 17740 88116 17746
rect 88064 17682 88116 17688
rect 88260 17134 88288 19774
rect 88352 19774 88426 19802
rect 88536 19774 88610 19802
rect 88720 19774 88794 19802
rect 88904 19774 88978 19802
rect 89088 19774 89162 19802
rect 89272 19774 89346 19802
rect 89456 19774 89530 19802
rect 89640 19774 89714 19802
rect 89824 19774 89898 19802
rect 90008 19774 90082 19802
rect 90192 19774 90266 19802
rect 90376 19774 90450 19802
rect 90560 19774 90634 19802
rect 90790 19802 90818 20060
rect 90974 19802 91002 20060
rect 91158 19802 91186 20060
rect 91342 19802 91370 20060
rect 91526 19802 91554 20060
rect 91710 19802 91738 20060
rect 91894 19802 91922 20060
rect 92078 19802 92106 20060
rect 92262 19802 92290 20060
rect 92446 19802 92474 20060
rect 92630 19802 92658 20060
rect 90790 19774 90864 19802
rect 90974 19774 91048 19802
rect 91158 19774 91232 19802
rect 88248 17128 88300 17134
rect 88248 17070 88300 17076
rect 87788 15224 87840 15230
rect 87788 15166 87840 15172
rect 88248 14272 88300 14278
rect 88248 14214 88300 14220
rect 87972 12844 88024 12850
rect 87972 12786 88024 12792
rect 87984 9246 88012 12786
rect 88260 9926 88288 14214
rect 88352 10588 88380 19774
rect 88536 11830 88564 19774
rect 88524 11824 88576 11830
rect 88524 11766 88576 11772
rect 88352 10560 88564 10588
rect 88340 10328 88392 10334
rect 88340 10270 88392 10276
rect 88430 10296 88486 10305
rect 88248 9920 88300 9926
rect 88248 9862 88300 9868
rect 87972 9240 88024 9246
rect 87972 9182 88024 9188
rect 88352 9110 88380 10270
rect 88430 10231 88486 10240
rect 88340 9104 88392 9110
rect 88340 9046 88392 9052
rect 88444 8945 88472 10231
rect 88430 8936 88486 8945
rect 88430 8871 88486 8880
rect 88432 8696 88484 8702
rect 88432 8638 88484 8644
rect 88340 6724 88392 6730
rect 88340 6666 88392 6672
rect 87696 6180 87748 6186
rect 87696 6122 87748 6128
rect 87972 4888 88024 4894
rect 87972 4830 88024 4836
rect 87604 2304 87656 2310
rect 87604 2246 87656 2252
rect 87144 2236 87196 2242
rect 87144 2178 87196 2184
rect 87156 814 87184 2178
rect 87144 808 87196 814
rect 87144 750 87196 756
rect 87984 480 88012 4830
rect 88352 4049 88380 6666
rect 88338 4040 88394 4049
rect 88338 3975 88394 3984
rect 88444 3534 88472 8638
rect 88536 5030 88564 10560
rect 88720 7682 88748 19774
rect 88800 17196 88852 17202
rect 88800 17138 88852 17144
rect 88812 12034 88840 17138
rect 88904 12034 88932 19774
rect 88984 15224 89036 15230
rect 88984 15166 89036 15172
rect 88800 12028 88852 12034
rect 88800 11970 88852 11976
rect 88892 12028 88944 12034
rect 88892 11970 88944 11976
rect 88996 10810 89024 15166
rect 89088 14550 89116 19774
rect 89272 17542 89300 19774
rect 89260 17536 89312 17542
rect 89260 17478 89312 17484
rect 89456 16182 89484 19774
rect 89534 17232 89590 17241
rect 89534 17167 89590 17176
rect 89548 16425 89576 17167
rect 89534 16416 89590 16425
rect 89534 16351 89590 16360
rect 89444 16176 89496 16182
rect 89444 16118 89496 16124
rect 89640 15450 89668 19774
rect 89720 17808 89772 17814
rect 89720 17750 89772 17756
rect 89548 15422 89668 15450
rect 89076 14544 89128 14550
rect 89076 14486 89128 14492
rect 89548 12510 89576 15422
rect 89628 15292 89680 15298
rect 89628 15234 89680 15240
rect 89640 14906 89668 15234
rect 89732 15026 89760 17750
rect 89720 15020 89772 15026
rect 89720 14962 89772 14968
rect 89640 14878 89760 14906
rect 89536 12504 89588 12510
rect 89536 12446 89588 12452
rect 88984 10804 89036 10810
rect 88984 10746 89036 10752
rect 88708 7676 88760 7682
rect 88708 7618 88760 7624
rect 88616 6656 88668 6662
rect 88616 6598 88668 6604
rect 88628 5982 88656 6598
rect 88616 5976 88668 5982
rect 88616 5918 88668 5924
rect 88524 5024 88576 5030
rect 88524 4966 88576 4972
rect 89168 3732 89220 3738
rect 89168 3674 89220 3680
rect 88432 3528 88484 3534
rect 88432 3470 88484 3476
rect 89180 480 89208 3674
rect 79324 128 79376 134
rect 79324 70 79376 76
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89732 354 89760 14878
rect 89824 1193 89852 19774
rect 89904 15632 89956 15638
rect 89904 15574 89956 15580
rect 89916 13462 89944 15574
rect 89904 13456 89956 13462
rect 89904 13398 89956 13404
rect 90008 5982 90036 19774
rect 90088 17604 90140 17610
rect 90088 17546 90140 17552
rect 90100 10606 90128 17546
rect 90192 16574 90220 19774
rect 90376 17950 90404 19774
rect 90364 17944 90416 17950
rect 90364 17886 90416 17892
rect 90192 16546 90312 16574
rect 90180 15224 90232 15230
rect 90180 15166 90232 15172
rect 90088 10600 90140 10606
rect 90088 10542 90140 10548
rect 90192 9450 90220 15166
rect 90180 9444 90232 9450
rect 90180 9386 90232 9392
rect 90180 7812 90232 7818
rect 90180 7754 90232 7760
rect 89996 5976 90048 5982
rect 89996 5918 90048 5924
rect 90192 3874 90220 7754
rect 90284 7750 90312 16546
rect 90364 15700 90416 15706
rect 90364 15642 90416 15648
rect 90376 8022 90404 15642
rect 90560 14958 90588 19774
rect 90732 17400 90784 17406
rect 90732 17342 90784 17348
rect 90744 16289 90772 17342
rect 90730 16280 90786 16289
rect 90836 16250 90864 19774
rect 91020 16998 91048 19774
rect 91008 16992 91060 16998
rect 91008 16934 91060 16940
rect 91204 16930 91232 19774
rect 91296 19774 91370 19802
rect 91480 19774 91554 19802
rect 91664 19774 91738 19802
rect 91848 19774 91922 19802
rect 92032 19774 92106 19802
rect 92216 19774 92290 19802
rect 92400 19774 92474 19802
rect 92584 19774 92658 19802
rect 92814 19802 92842 20060
rect 92998 19802 93026 20060
rect 93182 19802 93210 20060
rect 92814 19774 92888 19802
rect 91192 16924 91244 16930
rect 91192 16866 91244 16872
rect 91008 16856 91060 16862
rect 91008 16798 91060 16804
rect 90730 16215 90786 16224
rect 90824 16244 90876 16250
rect 90824 16186 90876 16192
rect 91020 15774 91048 16798
rect 91296 16114 91324 19774
rect 91374 18048 91430 18057
rect 91374 17983 91430 17992
rect 91388 17202 91416 17983
rect 91480 17814 91508 19774
rect 91468 17808 91520 17814
rect 91468 17750 91520 17756
rect 91560 17740 91612 17746
rect 91560 17682 91612 17688
rect 91376 17196 91428 17202
rect 91376 17138 91428 17144
rect 91284 16108 91336 16114
rect 91284 16050 91336 16056
rect 91008 15768 91060 15774
rect 91008 15710 91060 15716
rect 90548 14952 90600 14958
rect 90548 14894 90600 14900
rect 91098 14920 91154 14929
rect 91098 14855 91154 14864
rect 91112 12646 91140 14855
rect 91572 13258 91600 17682
rect 91560 13252 91612 13258
rect 91560 13194 91612 13200
rect 91664 13190 91692 19774
rect 91744 16856 91796 16862
rect 91744 16798 91796 16804
rect 91756 16386 91784 16798
rect 91744 16380 91796 16386
rect 91744 16322 91796 16328
rect 91744 15836 91796 15842
rect 91744 15778 91796 15784
rect 91652 13184 91704 13190
rect 91652 13126 91704 13132
rect 91192 12980 91244 12986
rect 91192 12922 91244 12928
rect 91100 12640 91152 12646
rect 91100 12582 91152 12588
rect 90640 12504 90692 12510
rect 90640 12446 90692 12452
rect 90364 8016 90416 8022
rect 90364 7958 90416 7964
rect 90652 7818 90680 12446
rect 91008 9716 91060 9722
rect 91008 9658 91060 9664
rect 91020 9586 91048 9658
rect 91008 9580 91060 9586
rect 91008 9522 91060 9528
rect 91204 9353 91232 12922
rect 91652 9648 91704 9654
rect 91652 9590 91704 9596
rect 91190 9344 91246 9353
rect 91190 9279 91246 9288
rect 91008 8968 91060 8974
rect 91008 8910 91060 8916
rect 91020 8702 91048 8910
rect 91008 8696 91060 8702
rect 91008 8638 91060 8644
rect 90640 7812 90692 7818
rect 90640 7754 90692 7760
rect 90272 7744 90324 7750
rect 90272 7686 90324 7692
rect 90180 3868 90232 3874
rect 90180 3810 90232 3816
rect 91560 3324 91612 3330
rect 91560 3266 91612 3272
rect 89810 1184 89866 1193
rect 89810 1119 89866 1128
rect 91572 480 91600 3266
rect 91664 2242 91692 9590
rect 91756 3126 91784 15778
rect 91848 9450 91876 19774
rect 92032 15842 92060 19774
rect 92020 15836 92072 15842
rect 92020 15778 92072 15784
rect 91836 9444 91888 9450
rect 91836 9386 91888 9392
rect 92216 6390 92244 19774
rect 92400 18306 92428 19774
rect 92308 18278 92428 18306
rect 92308 10470 92336 18278
rect 92584 17898 92612 19774
rect 92400 17870 92612 17898
rect 92400 13938 92428 17870
rect 92572 17808 92624 17814
rect 92572 17750 92624 17756
rect 92584 15230 92612 17750
rect 92860 17542 92888 19774
rect 92952 19774 93026 19802
rect 93136 19774 93210 19802
rect 93366 19802 93394 20060
rect 93550 19802 93578 20060
rect 93734 19802 93762 20060
rect 93918 19802 93946 20060
rect 93366 19774 93440 19802
rect 92848 17536 92900 17542
rect 92848 17478 92900 17484
rect 92572 15224 92624 15230
rect 92572 15166 92624 15172
rect 92756 15224 92808 15230
rect 92756 15166 92808 15172
rect 92570 14648 92626 14657
rect 92570 14583 92626 14592
rect 92388 13932 92440 13938
rect 92388 13874 92440 13880
rect 92584 11665 92612 14583
rect 92570 11656 92626 11665
rect 92570 11591 92626 11600
rect 92296 10464 92348 10470
rect 92296 10406 92348 10412
rect 92480 10124 92532 10130
rect 92480 10066 92532 10072
rect 92204 6384 92256 6390
rect 92204 6326 92256 6332
rect 92388 6316 92440 6322
rect 92388 6258 92440 6264
rect 92400 3194 92428 6258
rect 92492 3738 92520 10066
rect 92768 7886 92796 15166
rect 92952 11082 92980 19774
rect 93136 17814 93164 19774
rect 93124 17808 93176 17814
rect 93124 17750 93176 17756
rect 93124 17672 93176 17678
rect 93124 17614 93176 17620
rect 92940 11076 92992 11082
rect 92940 11018 92992 11024
rect 92756 7880 92808 7886
rect 92756 7822 92808 7828
rect 92572 6384 92624 6390
rect 92572 6326 92624 6332
rect 92584 5982 92612 6326
rect 92572 5976 92624 5982
rect 92572 5918 92624 5924
rect 92756 3868 92808 3874
rect 92756 3810 92808 3816
rect 92480 3732 92532 3738
rect 92480 3674 92532 3680
rect 92388 3188 92440 3194
rect 92388 3130 92440 3136
rect 91744 3120 91796 3126
rect 91744 3062 91796 3068
rect 91652 2236 91704 2242
rect 91652 2178 91704 2184
rect 92768 480 92796 3810
rect 92940 3664 92992 3670
rect 92940 3606 92992 3612
rect 92952 3330 92980 3606
rect 92940 3324 92992 3330
rect 92940 3266 92992 3272
rect 93136 2145 93164 17614
rect 93412 16726 93440 19774
rect 93504 19774 93578 19802
rect 93688 19774 93762 19802
rect 93872 19774 93946 19802
rect 94102 19802 94130 20060
rect 94286 19802 94314 20060
rect 94470 19802 94498 20060
rect 94654 19802 94682 20060
rect 94838 19802 94866 20060
rect 95022 19802 95050 20060
rect 95206 19938 95234 20060
rect 94102 19774 94176 19802
rect 93400 16720 93452 16726
rect 93400 16662 93452 16668
rect 93504 14142 93532 19774
rect 93584 16924 93636 16930
rect 93584 16866 93636 16872
rect 93596 14278 93624 16866
rect 93584 14272 93636 14278
rect 93584 14214 93636 14220
rect 93492 14136 93544 14142
rect 93492 14078 93544 14084
rect 93584 12028 93636 12034
rect 93584 11970 93636 11976
rect 93596 7274 93624 11970
rect 93584 7268 93636 7274
rect 93584 7210 93636 7216
rect 93122 2136 93178 2145
rect 93122 2071 93178 2080
rect 90334 354 90446 480
rect 89732 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93688 241 93716 19774
rect 93768 17128 93820 17134
rect 93768 17070 93820 17076
rect 93780 16930 93808 17070
rect 93768 16924 93820 16930
rect 93768 16866 93820 16872
rect 93872 16574 93900 19774
rect 94148 17610 94176 19774
rect 94240 19774 94314 19802
rect 94424 19774 94498 19802
rect 94608 19774 94682 19802
rect 94792 19774 94866 19802
rect 94976 19774 95050 19802
rect 95160 19910 95234 19938
rect 94240 19378 94268 19774
rect 94228 19372 94280 19378
rect 94228 19314 94280 19320
rect 94136 17604 94188 17610
rect 94136 17546 94188 17552
rect 94136 17468 94188 17474
rect 94136 17410 94188 17416
rect 93872 16546 93992 16574
rect 93964 12434 93992 16546
rect 94148 14929 94176 17410
rect 94134 14920 94190 14929
rect 94134 14855 94190 14864
rect 94424 13841 94452 19774
rect 94608 17950 94636 19774
rect 94596 17944 94648 17950
rect 94596 17886 94648 17892
rect 94688 16720 94740 16726
rect 94688 16662 94740 16668
rect 94594 15192 94650 15201
rect 94594 15127 94650 15136
rect 94410 13832 94466 13841
rect 94410 13767 94466 13776
rect 93964 12406 94084 12434
rect 93768 11756 93820 11762
rect 93768 11698 93820 11704
rect 93780 10130 93808 11698
rect 93768 10124 93820 10130
rect 93768 10066 93820 10072
rect 93860 9172 93912 9178
rect 93860 9114 93912 9120
rect 93872 3874 93900 9114
rect 94056 8090 94084 12406
rect 94504 10668 94556 10674
rect 94504 10610 94556 10616
rect 94516 10334 94544 10610
rect 94504 10328 94556 10334
rect 94504 10270 94556 10276
rect 94504 8696 94556 8702
rect 94504 8638 94556 8644
rect 94044 8084 94096 8090
rect 94044 8026 94096 8032
rect 94516 8022 94544 8638
rect 94608 8294 94636 15127
rect 94700 12034 94728 16662
rect 94688 12028 94740 12034
rect 94688 11970 94740 11976
rect 94792 9314 94820 19774
rect 94976 16574 95004 19774
rect 95160 18306 95188 19910
rect 95240 19848 95292 19854
rect 95240 19790 95292 19796
rect 95390 19802 95418 20060
rect 95574 19802 95602 20060
rect 95758 19802 95786 20060
rect 95942 19854 95970 20060
rect 95068 18278 95188 18306
rect 95068 17202 95096 18278
rect 95148 18216 95200 18222
rect 95148 18158 95200 18164
rect 95056 17196 95108 17202
rect 95056 17138 95108 17144
rect 95160 17066 95188 18158
rect 95148 17060 95200 17066
rect 95148 17002 95200 17008
rect 94976 16546 95096 16574
rect 94962 15328 95018 15337
rect 94962 15263 95018 15272
rect 94976 12345 95004 15263
rect 94962 12336 95018 12345
rect 94962 12271 95018 12280
rect 95068 11490 95096 16546
rect 95146 14784 95202 14793
rect 95146 14719 95202 14728
rect 95160 12481 95188 14719
rect 95146 12472 95202 12481
rect 95146 12407 95202 12416
rect 95252 12434 95280 19790
rect 95390 19774 95464 19802
rect 95252 12406 95372 12434
rect 95238 11928 95294 11937
rect 95238 11863 95294 11872
rect 95056 11484 95108 11490
rect 95056 11426 95108 11432
rect 95056 11076 95108 11082
rect 95056 11018 95108 11024
rect 94780 9308 94832 9314
rect 94780 9250 94832 9256
rect 94596 8288 94648 8294
rect 94596 8230 94648 8236
rect 94504 8016 94556 8022
rect 94504 7958 94556 7964
rect 94504 7676 94556 7682
rect 94504 7618 94556 7624
rect 94516 5914 94544 7618
rect 94504 5908 94556 5914
rect 94504 5850 94556 5856
rect 95068 5409 95096 11018
rect 95252 10305 95280 11863
rect 95238 10296 95294 10305
rect 95238 10231 95294 10240
rect 95240 9036 95292 9042
rect 95240 8978 95292 8984
rect 95252 7206 95280 8978
rect 95344 8498 95372 12406
rect 95436 11082 95464 19774
rect 95528 19774 95602 19802
rect 95712 19774 95786 19802
rect 95930 19848 95982 19854
rect 96126 19802 96154 20060
rect 96310 19802 96338 20060
rect 96494 19802 96522 20060
rect 96678 19802 96706 20060
rect 96862 19938 96890 20060
rect 95930 19790 95982 19796
rect 96080 19774 96154 19802
rect 96264 19774 96338 19802
rect 96448 19774 96522 19802
rect 96632 19774 96706 19802
rect 96816 19910 96890 19938
rect 95528 16386 95556 19774
rect 95712 17134 95740 19774
rect 95790 17232 95846 17241
rect 95790 17167 95846 17176
rect 95700 17128 95752 17134
rect 95700 17070 95752 17076
rect 95516 16380 95568 16386
rect 95516 16322 95568 16328
rect 95804 15230 95832 17167
rect 95792 15224 95844 15230
rect 95792 15166 95844 15172
rect 95790 13560 95846 13569
rect 95790 13495 95846 13504
rect 95424 11076 95476 11082
rect 95424 11018 95476 11024
rect 95804 10849 95832 13495
rect 95790 10840 95846 10849
rect 95790 10775 95846 10784
rect 95424 10668 95476 10674
rect 95424 10610 95476 10616
rect 95332 8492 95384 8498
rect 95332 8434 95384 8440
rect 95240 7200 95292 7206
rect 95240 7142 95292 7148
rect 95436 6866 95464 10610
rect 96080 8294 96108 19774
rect 96068 8288 96120 8294
rect 96068 8230 96120 8236
rect 95424 6860 95476 6866
rect 95424 6802 95476 6808
rect 96264 6769 96292 19774
rect 96342 14784 96398 14793
rect 96342 14719 96398 14728
rect 96356 13705 96384 14719
rect 96342 13696 96398 13705
rect 96342 13631 96398 13640
rect 96448 12442 96476 19774
rect 96528 19372 96580 19378
rect 96528 19314 96580 19320
rect 96540 19281 96568 19314
rect 96526 19272 96582 19281
rect 96526 19207 96582 19216
rect 96526 14512 96582 14521
rect 96526 14447 96582 14456
rect 96540 13705 96568 14447
rect 96526 13696 96582 13705
rect 96526 13631 96582 13640
rect 96526 13016 96582 13025
rect 96526 12951 96582 12960
rect 96436 12436 96488 12442
rect 96436 12378 96488 12384
rect 96540 12209 96568 12951
rect 96632 12434 96660 19774
rect 96712 17944 96764 17950
rect 96712 17886 96764 17892
rect 96724 16862 96752 17886
rect 96712 16856 96764 16862
rect 96712 16798 96764 16804
rect 96632 12406 96752 12434
rect 96526 12200 96582 12209
rect 96526 12135 96582 12144
rect 96620 10532 96672 10538
rect 96620 10474 96672 10480
rect 96632 10334 96660 10474
rect 96344 10328 96396 10334
rect 96344 10270 96396 10276
rect 96620 10328 96672 10334
rect 96620 10270 96672 10276
rect 96250 6760 96306 6769
rect 96250 6695 96306 6704
rect 95238 6216 95294 6225
rect 95238 6151 95294 6160
rect 95054 5400 95110 5409
rect 95054 5335 95110 5344
rect 93860 3868 93912 3874
rect 93860 3810 93912 3816
rect 93952 3732 94004 3738
rect 93952 3674 94004 3680
rect 93964 480 93992 3674
rect 95148 3256 95200 3262
rect 95148 3198 95200 3204
rect 95160 480 95188 3198
rect 95252 2825 95280 6151
rect 96356 3670 96384 10270
rect 96620 8696 96672 8702
rect 96620 8638 96672 8644
rect 96632 7138 96660 8638
rect 96724 7682 96752 12406
rect 96816 10674 96844 19910
rect 97046 19802 97074 20060
rect 97230 19802 97258 20060
rect 97414 19802 97442 20060
rect 97598 19802 97626 20060
rect 97782 19802 97810 20060
rect 97966 19938 97994 20060
rect 96908 19774 97074 19802
rect 97184 19774 97258 19802
rect 97368 19774 97442 19802
rect 97552 19774 97626 19802
rect 97736 19774 97810 19802
rect 97920 19910 97994 19938
rect 96908 16454 96936 19774
rect 97080 17604 97132 17610
rect 97080 17546 97132 17552
rect 96896 16448 96948 16454
rect 96896 16390 96948 16396
rect 97092 14521 97120 17546
rect 97184 14657 97212 19774
rect 97368 17785 97396 19774
rect 97354 17776 97410 17785
rect 97354 17711 97410 17720
rect 97264 17604 97316 17610
rect 97264 17546 97316 17552
rect 97276 17406 97304 17546
rect 97552 17474 97580 19774
rect 97540 17468 97592 17474
rect 97540 17410 97592 17416
rect 97264 17400 97316 17406
rect 97264 17342 97316 17348
rect 97356 17400 97408 17406
rect 97356 17342 97408 17348
rect 97264 16040 97316 16046
rect 97264 15982 97316 15988
rect 97170 14648 97226 14657
rect 97170 14583 97226 14592
rect 97078 14512 97134 14521
rect 97078 14447 97134 14456
rect 96894 13832 96950 13841
rect 96894 13767 96950 13776
rect 96908 11014 96936 13767
rect 96896 11008 96948 11014
rect 96896 10950 96948 10956
rect 96804 10668 96856 10674
rect 96804 10610 96856 10616
rect 96804 10532 96856 10538
rect 96804 10474 96856 10480
rect 96712 7676 96764 7682
rect 96712 7618 96764 7624
rect 96620 7132 96672 7138
rect 96620 7074 96672 7080
rect 96816 6633 96844 10474
rect 96896 10328 96948 10334
rect 96896 10270 96948 10276
rect 96802 6624 96858 6633
rect 96802 6559 96858 6568
rect 96344 3664 96396 3670
rect 96344 3606 96396 3612
rect 96908 3602 96936 10270
rect 96896 3596 96948 3602
rect 96896 3538 96948 3544
rect 97276 3330 97304 15982
rect 97368 5506 97396 17342
rect 97632 16720 97684 16726
rect 97632 16662 97684 16668
rect 97540 14272 97592 14278
rect 97540 14214 97592 14220
rect 97552 11234 97580 14214
rect 97644 12434 97672 16662
rect 97736 15638 97764 19774
rect 97814 18184 97870 18193
rect 97814 18119 97870 18128
rect 97828 16998 97856 18119
rect 97920 17950 97948 19910
rect 98150 19802 98178 20060
rect 98334 19802 98362 20060
rect 98518 19802 98546 20060
rect 98702 19802 98730 20060
rect 98886 19802 98914 20060
rect 99070 19802 99098 20060
rect 99254 19802 99282 20060
rect 99438 19802 99466 20060
rect 99622 19802 99650 20060
rect 99806 19802 99834 20060
rect 98012 19774 98178 19802
rect 98288 19774 98362 19802
rect 98472 19774 98546 19802
rect 98656 19774 98730 19802
rect 98840 19774 98914 19802
rect 99024 19774 99098 19802
rect 99208 19774 99282 19802
rect 99392 19774 99466 19802
rect 99576 19774 99650 19802
rect 99760 19774 99834 19802
rect 99990 19802 100018 20060
rect 100174 19802 100202 20060
rect 100358 19802 100386 20060
rect 100542 19802 100570 20060
rect 100726 19802 100754 20060
rect 100910 19938 100938 20060
rect 99990 19774 100064 19802
rect 97908 17944 97960 17950
rect 97908 17886 97960 17892
rect 97908 17740 97960 17746
rect 97908 17682 97960 17688
rect 97816 16992 97868 16998
rect 97816 16934 97868 16940
rect 97816 16856 97868 16862
rect 97816 16798 97868 16804
rect 97724 15632 97776 15638
rect 97724 15574 97776 15580
rect 97828 13569 97856 16798
rect 97920 16658 97948 17682
rect 97908 16652 97960 16658
rect 97908 16594 97960 16600
rect 98012 15450 98040 19774
rect 98092 18284 98144 18290
rect 98092 18226 98144 18232
rect 98104 15706 98132 18226
rect 98288 16046 98316 19774
rect 98276 16040 98328 16046
rect 98276 15982 98328 15988
rect 98276 15836 98328 15842
rect 98276 15778 98328 15784
rect 98092 15700 98144 15706
rect 98092 15642 98144 15648
rect 98184 15632 98236 15638
rect 98184 15574 98236 15580
rect 98012 15422 98132 15450
rect 97814 13560 97870 13569
rect 97814 13495 97870 13504
rect 97644 12406 97764 12434
rect 97552 11206 97672 11234
rect 97540 11076 97592 11082
rect 97540 11018 97592 11024
rect 97448 8288 97500 8294
rect 97448 8230 97500 8236
rect 97460 6254 97488 8230
rect 97448 6248 97500 6254
rect 97448 6190 97500 6196
rect 97356 5500 97408 5506
rect 97356 5442 97408 5448
rect 97448 3868 97500 3874
rect 97448 3810 97500 3816
rect 96252 3324 96304 3330
rect 96252 3266 96304 3272
rect 97264 3324 97316 3330
rect 97264 3266 97316 3272
rect 95238 2816 95294 2825
rect 95238 2751 95294 2760
rect 96264 480 96292 3266
rect 97460 480 97488 3810
rect 97552 1902 97580 11018
rect 97644 5545 97672 11206
rect 97736 9042 97764 12406
rect 98104 10985 98132 15422
rect 98196 13297 98224 15574
rect 98182 13288 98238 13297
rect 98182 13223 98238 13232
rect 98090 10976 98146 10985
rect 98090 10911 98146 10920
rect 98092 10124 98144 10130
rect 98092 10066 98144 10072
rect 98000 9172 98052 9178
rect 98000 9114 98052 9120
rect 97724 9036 97776 9042
rect 97724 8978 97776 8984
rect 98012 8129 98040 9114
rect 98104 8294 98132 10066
rect 98288 9654 98316 15778
rect 98276 9648 98328 9654
rect 98276 9590 98328 9596
rect 98092 8288 98144 8294
rect 98092 8230 98144 8236
rect 97998 8120 98054 8129
rect 97998 8055 98054 8064
rect 97998 7576 98054 7585
rect 97998 7511 98054 7520
rect 98012 6905 98040 7511
rect 97998 6896 98054 6905
rect 97998 6831 98054 6840
rect 98472 6633 98500 19774
rect 98656 10334 98684 19774
rect 98736 17944 98788 17950
rect 98736 17886 98788 17892
rect 98644 10328 98696 10334
rect 98644 10270 98696 10276
rect 98748 9489 98776 17886
rect 98734 9480 98790 9489
rect 98734 9415 98790 9424
rect 98458 6624 98514 6633
rect 98458 6559 98514 6568
rect 98840 6497 98868 19774
rect 99024 18290 99052 19774
rect 99208 19446 99236 19774
rect 99196 19440 99248 19446
rect 99196 19382 99248 19388
rect 99012 18284 99064 18290
rect 99012 18226 99064 18232
rect 99288 17536 99340 17542
rect 99288 17478 99340 17484
rect 99196 17332 99248 17338
rect 99196 17274 99248 17280
rect 99208 15706 99236 17274
rect 99300 16454 99328 17478
rect 99288 16448 99340 16454
rect 99288 16390 99340 16396
rect 99196 15700 99248 15706
rect 99196 15642 99248 15648
rect 99392 15230 99420 19774
rect 99472 17672 99524 17678
rect 99472 17614 99524 17620
rect 99484 15337 99512 17614
rect 99470 15328 99526 15337
rect 99470 15263 99526 15272
rect 99380 15224 99432 15230
rect 99380 15166 99432 15172
rect 98826 6488 98882 6497
rect 98826 6423 98882 6432
rect 98000 5908 98052 5914
rect 98000 5850 98052 5856
rect 97630 5536 97686 5545
rect 97630 5471 97686 5480
rect 98012 3262 98040 5850
rect 98644 3392 98696 3398
rect 99576 3369 99604 19774
rect 98644 3334 98696 3340
rect 99562 3360 99618 3369
rect 98000 3256 98052 3262
rect 98000 3198 98052 3204
rect 97540 1896 97592 1902
rect 97540 1838 97592 1844
rect 98656 480 98684 3334
rect 99562 3295 99618 3304
rect 99760 921 99788 19774
rect 100036 17338 100064 19774
rect 100128 19774 100202 19802
rect 100312 19774 100386 19802
rect 100496 19774 100570 19802
rect 100680 19774 100754 19802
rect 100864 19910 100938 19938
rect 100128 17950 100156 19774
rect 100116 17944 100168 17950
rect 100116 17886 100168 17892
rect 100024 17332 100076 17338
rect 100024 17274 100076 17280
rect 100312 10577 100340 19774
rect 100298 10568 100354 10577
rect 100298 10503 100354 10512
rect 100392 9648 100444 9654
rect 100392 9590 100444 9596
rect 99840 3392 99892 3398
rect 99840 3334 99892 3340
rect 99746 912 99802 921
rect 99746 847 99802 856
rect 99852 480 99880 3334
rect 100404 2009 100432 9590
rect 100496 5273 100524 19774
rect 100680 18306 100708 19774
rect 100864 18494 100892 19910
rect 100944 19848 100996 19854
rect 101094 19802 101122 20060
rect 101278 19802 101306 20060
rect 101462 19802 101490 20060
rect 101646 19802 101674 20060
rect 101830 19802 101858 20060
rect 102014 19854 102042 20060
rect 100944 19790 100996 19796
rect 100852 18488 100904 18494
rect 100852 18430 100904 18436
rect 100588 18278 100708 18306
rect 100852 18284 100904 18290
rect 100588 15881 100616 18278
rect 100852 18226 100904 18232
rect 100758 18048 100814 18057
rect 100758 17983 100814 17992
rect 100772 16998 100800 17983
rect 100760 16992 100812 16998
rect 100760 16934 100812 16940
rect 100574 15872 100630 15881
rect 100574 15807 100630 15816
rect 100864 12209 100892 18226
rect 100850 12200 100906 12209
rect 100850 12135 100906 12144
rect 100760 11008 100812 11014
rect 100760 10950 100812 10956
rect 100772 9110 100800 10950
rect 100760 9104 100812 9110
rect 100760 9046 100812 9052
rect 100956 8702 100984 19790
rect 101048 19774 101122 19802
rect 101232 19774 101306 19802
rect 101416 19774 101490 19802
rect 101600 19774 101674 19802
rect 101784 19774 101858 19802
rect 102002 19848 102054 19854
rect 102002 19790 102054 19796
rect 102198 19802 102226 20060
rect 102382 19938 102410 20060
rect 102336 19910 102410 19938
rect 102566 19938 102594 20060
rect 102566 19910 102640 19938
rect 102198 19774 102272 19802
rect 101048 9654 101076 19774
rect 101128 18964 101180 18970
rect 101128 18906 101180 18912
rect 101140 17610 101168 18906
rect 101128 17604 101180 17610
rect 101128 17546 101180 17552
rect 101232 15337 101260 19774
rect 101312 18488 101364 18494
rect 101312 18430 101364 18436
rect 101324 16862 101352 18430
rect 101416 18290 101444 19774
rect 101404 18284 101456 18290
rect 101404 18226 101456 18232
rect 101496 17196 101548 17202
rect 101496 17138 101548 17144
rect 101312 16856 101364 16862
rect 101312 16798 101364 16804
rect 101218 15328 101274 15337
rect 101218 15263 101274 15272
rect 101508 11937 101536 17138
rect 101600 16289 101628 19774
rect 101586 16280 101642 16289
rect 101586 16215 101642 16224
rect 101588 15224 101640 15230
rect 101588 15166 101640 15172
rect 101494 11928 101550 11937
rect 101494 11863 101550 11872
rect 101036 9648 101088 9654
rect 101036 9590 101088 9596
rect 101600 8974 101628 15166
rect 101680 10668 101732 10674
rect 101680 10610 101732 10616
rect 101220 8968 101272 8974
rect 101588 8968 101640 8974
rect 101220 8910 101272 8916
rect 101402 8936 101458 8945
rect 100944 8696 100996 8702
rect 100944 8638 100996 8644
rect 100482 5264 100538 5273
rect 100482 5199 100538 5208
rect 101232 3874 101260 8910
rect 101588 8910 101640 8916
rect 101402 8871 101458 8880
rect 101312 8764 101364 8770
rect 101312 8706 101364 8712
rect 101220 3868 101272 3874
rect 101220 3810 101272 3816
rect 101036 3800 101088 3806
rect 101036 3742 101088 3748
rect 100390 2000 100446 2009
rect 100390 1935 100446 1944
rect 100760 1964 100812 1970
rect 100760 1906 100812 1912
rect 100772 542 100800 1906
rect 100760 536 100812 542
rect 93674 232 93730 241
rect 93674 167 93730 176
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100760 478 100812 484
rect 101048 480 101076 3742
rect 101324 3262 101352 8706
rect 101416 6866 101444 8871
rect 101404 6860 101456 6866
rect 101404 6802 101456 6808
rect 101692 4554 101720 10610
rect 101680 4548 101732 4554
rect 101680 4490 101732 4496
rect 101784 4185 101812 19774
rect 102140 18284 102192 18290
rect 102140 18226 102192 18232
rect 102152 17882 102180 18226
rect 102140 17876 102192 17882
rect 102140 17818 102192 17824
rect 102244 17490 102272 19774
rect 102336 17678 102364 19910
rect 102612 19582 102640 19910
rect 102750 19802 102778 20060
rect 102934 19802 102962 20060
rect 103118 19802 103146 20060
rect 103302 19802 103330 20060
rect 103486 19802 103514 20060
rect 102704 19774 102778 19802
rect 102888 19774 102962 19802
rect 103072 19774 103146 19802
rect 103256 19774 103330 19802
rect 103440 19774 103514 19802
rect 103670 19802 103698 20060
rect 103854 19802 103882 20060
rect 104038 19802 104066 20060
rect 104222 19802 104250 20060
rect 104406 19802 104434 20060
rect 104590 19802 104618 20060
rect 104774 19802 104802 20060
rect 103670 19774 103744 19802
rect 102600 19576 102652 19582
rect 102600 19518 102652 19524
rect 102324 17672 102376 17678
rect 102324 17614 102376 17620
rect 102244 17462 102548 17490
rect 102324 17060 102376 17066
rect 102324 17002 102376 17008
rect 102140 13864 102192 13870
rect 102140 13806 102192 13812
rect 102152 12782 102180 13806
rect 102140 12776 102192 12782
rect 102140 12718 102192 12724
rect 102140 12504 102192 12510
rect 102140 12446 102192 12452
rect 102152 9586 102180 12446
rect 102336 10674 102364 17002
rect 102416 16856 102468 16862
rect 102416 16798 102468 16804
rect 102428 11801 102456 16798
rect 102414 11792 102470 11801
rect 102414 11727 102470 11736
rect 102324 10668 102376 10674
rect 102324 10610 102376 10616
rect 102520 10441 102548 17462
rect 102506 10432 102562 10441
rect 102506 10367 102562 10376
rect 102140 9580 102192 9586
rect 102140 9522 102192 9528
rect 102140 8356 102192 8362
rect 102140 8298 102192 8304
rect 102152 7993 102180 8298
rect 102704 8294 102732 19774
rect 102600 8288 102652 8294
rect 102600 8230 102652 8236
rect 102692 8288 102744 8294
rect 102692 8230 102744 8236
rect 102138 7984 102194 7993
rect 102138 7919 102194 7928
rect 102138 7032 102194 7041
rect 102138 6967 102194 6976
rect 102152 6089 102180 6967
rect 102138 6080 102194 6089
rect 102138 6015 102194 6024
rect 101770 4176 101826 4185
rect 101770 4111 101826 4120
rect 102232 3596 102284 3602
rect 102232 3538 102284 3544
rect 101312 3256 101364 3262
rect 101312 3198 101364 3204
rect 102244 480 102272 3538
rect 102612 3194 102640 8230
rect 102888 3602 102916 19774
rect 102968 19372 103020 19378
rect 102968 19314 103020 19320
rect 102980 15842 103008 19314
rect 103072 17542 103100 19774
rect 103060 17536 103112 17542
rect 103060 17478 103112 17484
rect 102968 15836 103020 15842
rect 102968 15778 103020 15784
rect 103256 6361 103284 19774
rect 103440 17542 103468 19774
rect 103716 19514 103744 19774
rect 103808 19774 103882 19802
rect 103992 19774 104066 19802
rect 104176 19774 104250 19802
rect 104360 19774 104434 19802
rect 104544 19774 104618 19802
rect 104728 19774 104802 19802
rect 104958 19802 104986 20060
rect 105142 19802 105170 20060
rect 105326 19802 105354 20060
rect 105510 19802 105538 20060
rect 104958 19774 105032 19802
rect 103704 19508 103756 19514
rect 103704 19450 103756 19456
rect 103428 17536 103480 17542
rect 103428 17478 103480 17484
rect 103612 17468 103664 17474
rect 103612 17410 103664 17416
rect 103624 10538 103652 17410
rect 103704 17264 103756 17270
rect 103704 17206 103756 17212
rect 103716 11558 103744 17206
rect 103808 15881 103836 19774
rect 103794 15872 103850 15881
rect 103794 15807 103850 15816
rect 103704 11552 103756 11558
rect 103704 11494 103756 11500
rect 103612 10532 103664 10538
rect 103612 10474 103664 10480
rect 103520 9036 103572 9042
rect 103520 8978 103572 8984
rect 103242 6352 103298 6361
rect 103242 6287 103298 6296
rect 103532 5506 103560 8978
rect 103520 5500 103572 5506
rect 103520 5442 103572 5448
rect 103518 4312 103574 4321
rect 103518 4247 103574 4256
rect 103532 4049 103560 4247
rect 103518 4040 103574 4049
rect 103518 3975 103574 3984
rect 103336 3732 103388 3738
rect 103336 3674 103388 3680
rect 103428 3732 103480 3738
rect 103428 3674 103480 3680
rect 102876 3596 102928 3602
rect 102876 3538 102928 3544
rect 102600 3188 102652 3194
rect 102600 3130 102652 3136
rect 103348 480 103376 3674
rect 103440 3602 103468 3674
rect 103428 3596 103480 3602
rect 103428 3538 103480 3544
rect 103992 3058 104020 19774
rect 104176 17270 104204 19774
rect 104256 17808 104308 17814
rect 104256 17750 104308 17756
rect 104164 17264 104216 17270
rect 104164 17206 104216 17212
rect 104162 12880 104218 12889
rect 104162 12815 104218 12824
rect 104176 5137 104204 12815
rect 104268 8265 104296 17750
rect 104360 9217 104388 19774
rect 104440 19712 104492 19718
rect 104440 19654 104492 19660
rect 104452 15065 104480 19654
rect 104544 17134 104572 19774
rect 104728 19666 104756 19774
rect 104636 19638 104756 19666
rect 104532 17128 104584 17134
rect 104532 17070 104584 17076
rect 104636 16726 104664 19638
rect 104808 19372 104860 19378
rect 104808 19314 104860 19320
rect 104820 18193 104848 19314
rect 105004 18494 105032 19774
rect 105096 19774 105170 19802
rect 105280 19774 105354 19802
rect 105464 19774 105538 19802
rect 105694 19802 105722 20060
rect 105878 19802 105906 20060
rect 106062 19802 106090 20060
rect 106246 19802 106274 20060
rect 106430 19802 106458 20060
rect 106614 19802 106642 20060
rect 105694 19774 105768 19802
rect 104992 18488 105044 18494
rect 104992 18430 105044 18436
rect 104806 18184 104862 18193
rect 104806 18119 104862 18128
rect 104624 16720 104676 16726
rect 104624 16662 104676 16668
rect 104438 15056 104494 15065
rect 104438 14991 104494 15000
rect 104806 14512 104862 14521
rect 104806 14447 104862 14456
rect 104530 10704 104586 10713
rect 104820 10674 104848 14447
rect 104530 10639 104586 10648
rect 104808 10668 104860 10674
rect 104346 9208 104402 9217
rect 104346 9143 104402 9152
rect 104254 8256 104310 8265
rect 104254 8191 104310 8200
rect 104544 6905 104572 10639
rect 104808 10610 104860 10616
rect 104806 10296 104862 10305
rect 104806 10231 104862 10240
rect 104820 10062 104848 10231
rect 104808 10056 104860 10062
rect 104808 9998 104860 10004
rect 104898 7712 104954 7721
rect 104898 7647 104954 7656
rect 104530 6896 104586 6905
rect 104912 6866 104940 7647
rect 104530 6831 104586 6840
rect 104900 6860 104952 6866
rect 104900 6802 104952 6808
rect 104162 5128 104218 5137
rect 104162 5063 104218 5072
rect 104438 4856 104494 4865
rect 104438 4791 104494 4800
rect 104256 3868 104308 3874
rect 104256 3810 104308 3816
rect 103980 3052 104032 3058
rect 103980 2994 104032 3000
rect 104268 2553 104296 3810
rect 104452 3233 104480 4791
rect 104532 3664 104584 3670
rect 104532 3606 104584 3612
rect 104438 3224 104494 3233
rect 104438 3159 104494 3168
rect 104254 2544 104310 2553
rect 104254 2479 104310 2488
rect 104544 480 104572 3606
rect 105096 3602 105124 19774
rect 105176 18488 105228 18494
rect 105176 18430 105228 18436
rect 105188 14929 105216 18430
rect 105174 14920 105230 14929
rect 105174 14855 105230 14864
rect 105084 3596 105136 3602
rect 105084 3538 105136 3544
rect 104808 3392 104860 3398
rect 104808 3334 104860 3340
rect 104820 1970 104848 3334
rect 104808 1964 104860 1970
rect 104808 1906 104860 1912
rect 105280 1057 105308 19774
rect 105358 18320 105414 18329
rect 105358 18255 105414 18264
rect 105372 17610 105400 18255
rect 105360 17604 105412 17610
rect 105360 17546 105412 17552
rect 105464 13025 105492 19774
rect 105740 17610 105768 19774
rect 105832 19774 105906 19802
rect 106016 19774 106090 19802
rect 106200 19774 106274 19802
rect 106384 19774 106458 19802
rect 106568 19774 106642 19802
rect 106798 19802 106826 20060
rect 106982 19802 107010 20060
rect 107166 19802 107194 20060
rect 106798 19774 106872 19802
rect 105728 17604 105780 17610
rect 105728 17546 105780 17552
rect 105832 13705 105860 19774
rect 105818 13696 105874 13705
rect 105818 13631 105874 13640
rect 105450 13016 105506 13025
rect 105450 12951 105506 12960
rect 105636 12504 105688 12510
rect 105636 12446 105688 12452
rect 105648 11257 105676 12446
rect 105634 11248 105690 11257
rect 105634 11183 105690 11192
rect 106016 8129 106044 19774
rect 106094 18048 106150 18057
rect 106094 17983 106150 17992
rect 106108 16930 106136 17983
rect 106096 16924 106148 16930
rect 106096 16866 106148 16872
rect 106094 11656 106150 11665
rect 106094 11591 106150 11600
rect 106108 9761 106136 11591
rect 106094 9752 106150 9761
rect 106094 9687 106150 9696
rect 106002 8120 106058 8129
rect 106002 8055 106058 8064
rect 106200 3641 106228 19774
rect 106384 12442 106412 19774
rect 106372 12436 106424 12442
rect 106372 12378 106424 12384
rect 106280 11008 106332 11014
rect 106280 10950 106332 10956
rect 106292 9178 106320 10950
rect 106280 9172 106332 9178
rect 106280 9114 106332 9120
rect 106568 7993 106596 19774
rect 106844 17542 106872 19774
rect 106936 19774 107010 19802
rect 107120 19774 107194 19802
rect 107350 19802 107378 20060
rect 107534 19802 107562 20060
rect 107718 19802 107746 20060
rect 107350 19774 107424 19802
rect 106832 17536 106884 17542
rect 106832 17478 106884 17484
rect 106936 16862 106964 19774
rect 106924 16856 106976 16862
rect 106924 16798 106976 16804
rect 107120 16153 107148 19774
rect 107396 17882 107424 19774
rect 107488 19774 107562 19802
rect 107672 19774 107746 19802
rect 107902 19802 107930 20060
rect 108086 19802 108114 20060
rect 108270 19802 108298 20060
rect 108454 19802 108482 20060
rect 108638 19802 108666 20060
rect 108822 19802 108850 20060
rect 109006 19802 109034 20060
rect 109190 19938 109218 20060
rect 107902 19774 107976 19802
rect 107384 17876 107436 17882
rect 107384 17818 107436 17824
rect 107382 16688 107438 16697
rect 107382 16623 107438 16632
rect 107106 16144 107162 16153
rect 107106 16079 107162 16088
rect 107016 11620 107068 11626
rect 107016 11562 107068 11568
rect 106554 7984 106610 7993
rect 106554 7919 106610 7928
rect 106924 4140 106976 4146
rect 106924 4082 106976 4088
rect 106186 3632 106242 3641
rect 106186 3567 106242 3576
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 105266 1048 105322 1057
rect 105266 983 105322 992
rect 105740 480 105768 3062
rect 106188 2032 106240 2038
rect 106188 1974 106240 1980
rect 106200 882 106228 1974
rect 106188 876 106240 882
rect 106188 818 106240 824
rect 106936 480 106964 4082
rect 107028 3670 107056 11562
rect 107396 10849 107424 16623
rect 107488 12073 107516 19774
rect 107568 15836 107620 15842
rect 107568 15778 107620 15784
rect 107580 15201 107608 15778
rect 107566 15192 107622 15201
rect 107566 15127 107622 15136
rect 107566 13424 107622 13433
rect 107566 13359 107622 13368
rect 107580 13161 107608 13359
rect 107566 13152 107622 13161
rect 107566 13087 107622 13096
rect 107474 12064 107530 12073
rect 107474 11999 107530 12008
rect 107566 11928 107622 11937
rect 107566 11863 107622 11872
rect 107382 10840 107438 10849
rect 107382 10775 107438 10784
rect 107580 9042 107608 11863
rect 107568 9036 107620 9042
rect 107568 8978 107620 8984
rect 107476 8356 107528 8362
rect 107476 8298 107528 8304
rect 107488 4706 107516 8298
rect 107566 7032 107622 7041
rect 107566 6967 107622 6976
rect 107580 6866 107608 6967
rect 107568 6860 107620 6866
rect 107568 6802 107620 6808
rect 107672 6225 107700 19774
rect 107750 18184 107806 18193
rect 107750 18119 107806 18128
rect 107764 17746 107792 18119
rect 107752 17740 107804 17746
rect 107752 17682 107804 17688
rect 107948 16726 107976 19774
rect 108040 19774 108114 19802
rect 108224 19774 108298 19802
rect 108408 19774 108482 19802
rect 108592 19774 108666 19802
rect 108776 19774 108850 19802
rect 108960 19774 109034 19802
rect 109144 19910 109218 19938
rect 107936 16720 107988 16726
rect 107936 16662 107988 16668
rect 108040 14226 108068 19774
rect 108118 16824 108174 16833
rect 108118 16759 108174 16768
rect 107856 14198 108068 14226
rect 107750 12336 107806 12345
rect 107750 12271 107806 12280
rect 107764 9586 107792 12271
rect 107856 11762 107884 14198
rect 108132 14056 108160 16759
rect 107948 14028 108160 14056
rect 107844 11756 107896 11762
rect 107844 11698 107896 11704
rect 107948 11014 107976 14028
rect 108120 13864 108172 13870
rect 108120 13806 108172 13812
rect 108132 12986 108160 13806
rect 108120 12980 108172 12986
rect 108120 12922 108172 12928
rect 107936 11008 107988 11014
rect 107936 10950 107988 10956
rect 107752 9580 107804 9586
rect 107752 9522 107804 9528
rect 108026 7304 108082 7313
rect 108026 7239 108082 7248
rect 107658 6216 107714 6225
rect 107658 6151 107714 6160
rect 107488 4678 107700 4706
rect 107016 3664 107068 3670
rect 107016 3606 107068 3612
rect 107672 2553 107700 4678
rect 108040 4321 108068 7239
rect 108224 5137 108252 19774
rect 108304 17944 108356 17950
rect 108304 17886 108356 17892
rect 108316 17066 108344 17886
rect 108408 17814 108436 19774
rect 108396 17808 108448 17814
rect 108396 17750 108448 17756
rect 108304 17060 108356 17066
rect 108304 17002 108356 17008
rect 108304 14340 108356 14346
rect 108304 14282 108356 14288
rect 108316 13870 108344 14282
rect 108488 14068 108540 14074
rect 108488 14010 108540 14016
rect 108304 13864 108356 13870
rect 108304 13806 108356 13812
rect 108396 11688 108448 11694
rect 108396 11630 108448 11636
rect 108304 10532 108356 10538
rect 108304 10474 108356 10480
rect 108316 10334 108344 10474
rect 108304 10328 108356 10334
rect 108304 10270 108356 10276
rect 108408 10146 108436 11630
rect 108316 10118 108436 10146
rect 108210 5128 108266 5137
rect 108210 5063 108266 5072
rect 108026 4312 108082 4321
rect 108026 4247 108082 4256
rect 108212 3800 108264 3806
rect 108212 3742 108264 3748
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 107658 2544 107714 2553
rect 107658 2479 107714 2488
rect 108132 480 108160 3470
rect 108224 3398 108252 3742
rect 108316 3534 108344 10118
rect 108500 6914 108528 14010
rect 108592 11801 108620 19774
rect 108776 16574 108804 19774
rect 108960 17746 108988 19774
rect 109144 17746 109172 19910
rect 109224 19848 109276 19854
rect 109224 19790 109276 19796
rect 109374 19802 109402 20060
rect 109558 19802 109586 20060
rect 109742 19802 109770 20060
rect 108948 17740 109000 17746
rect 108948 17682 109000 17688
rect 109132 17740 109184 17746
rect 109132 17682 109184 17688
rect 108776 16546 109080 16574
rect 108578 11792 108634 11801
rect 108578 11727 108634 11736
rect 109052 10305 109080 16546
rect 109132 10668 109184 10674
rect 109132 10610 109184 10616
rect 109038 10296 109094 10305
rect 109038 10231 109094 10240
rect 109144 9178 109172 10610
rect 109132 9172 109184 9178
rect 109132 9114 109184 9120
rect 108948 7336 109000 7342
rect 108948 7278 109000 7284
rect 108408 6905 108528 6914
rect 108394 6896 108528 6905
rect 108450 6886 108528 6896
rect 108394 6831 108450 6840
rect 108396 4820 108448 4826
rect 108396 4762 108448 4768
rect 108408 3874 108436 4762
rect 108396 3868 108448 3874
rect 108396 3810 108448 3816
rect 108580 3868 108632 3874
rect 108580 3810 108632 3816
rect 108488 3800 108540 3806
rect 108488 3742 108540 3748
rect 108500 3602 108528 3742
rect 108488 3596 108540 3602
rect 108488 3538 108540 3544
rect 108304 3528 108356 3534
rect 108304 3470 108356 3476
rect 108212 3392 108264 3398
rect 108212 3334 108264 3340
rect 108592 3058 108620 3810
rect 108960 3602 108988 7278
rect 109236 5506 109264 19790
rect 109374 19774 109448 19802
rect 109420 15842 109448 19774
rect 109512 19774 109586 19802
rect 109696 19774 109770 19802
rect 109926 19802 109954 20060
rect 110110 19802 110138 20060
rect 110294 19854 110322 20060
rect 110282 19848 110334 19854
rect 109926 19774 110000 19802
rect 110110 19774 110184 19802
rect 110478 19802 110506 20060
rect 110282 19790 110334 19796
rect 109408 15836 109460 15842
rect 109408 15778 109460 15784
rect 109224 5500 109276 5506
rect 109224 5442 109276 5448
rect 109512 4146 109540 19774
rect 109592 17876 109644 17882
rect 109592 17818 109644 17824
rect 109604 12434 109632 17818
rect 109696 17474 109724 19774
rect 109684 17468 109736 17474
rect 109684 17410 109736 17416
rect 109776 17332 109828 17338
rect 109776 17274 109828 17280
rect 109604 12406 109724 12434
rect 109696 4894 109724 12406
rect 109788 7614 109816 17274
rect 109972 15609 110000 19774
rect 110156 17474 110184 19774
rect 110432 19774 110506 19802
rect 110662 19802 110690 20060
rect 110846 19938 110874 20060
rect 110800 19910 110874 19938
rect 110662 19774 110736 19802
rect 110144 17468 110196 17474
rect 110144 17410 110196 17416
rect 110326 16824 110382 16833
rect 110326 16759 110382 16768
rect 109958 15600 110014 15609
rect 109958 15535 110014 15544
rect 110340 15337 110368 16759
rect 110326 15328 110382 15337
rect 110326 15263 110382 15272
rect 110432 11665 110460 19774
rect 110510 18184 110566 18193
rect 110510 18119 110566 18128
rect 110524 17882 110552 18119
rect 110512 17876 110564 17882
rect 110512 17818 110564 17824
rect 110418 11656 110474 11665
rect 110418 11591 110474 11600
rect 110420 11484 110472 11490
rect 110420 11426 110472 11432
rect 110432 10674 110460 11426
rect 110510 11248 110566 11257
rect 110510 11183 110566 11192
rect 110420 10668 110472 10674
rect 110420 10610 110472 10616
rect 110524 8401 110552 11183
rect 110602 9616 110658 9625
rect 110602 9551 110658 9560
rect 110510 8392 110566 8401
rect 110510 8327 110566 8336
rect 109776 7608 109828 7614
rect 109776 7550 109828 7556
rect 110616 6089 110644 9551
rect 110602 6080 110658 6089
rect 110602 6015 110658 6024
rect 109684 4888 109736 4894
rect 109684 4830 109736 4836
rect 109500 4140 109552 4146
rect 109500 4082 109552 4088
rect 108948 3596 109000 3602
rect 108948 3538 109000 3544
rect 109316 3528 109368 3534
rect 110708 3505 110736 19774
rect 110800 17066 110828 19910
rect 111030 19802 111058 20060
rect 111214 19802 111242 20060
rect 111398 19802 111426 20060
rect 111582 19802 111610 20060
rect 111766 19802 111794 20060
rect 111950 19938 111978 20060
rect 111030 19774 111104 19802
rect 111214 19774 111288 19802
rect 110788 17060 110840 17066
rect 110788 17002 110840 17008
rect 111076 16522 111104 19774
rect 111156 19712 111208 19718
rect 111156 19654 111208 19660
rect 111064 16516 111116 16522
rect 111064 16458 111116 16464
rect 111064 15904 111116 15910
rect 111064 15846 111116 15852
rect 111076 3602 111104 15846
rect 111168 15065 111196 19654
rect 111260 16794 111288 19774
rect 111352 19774 111426 19802
rect 111536 19774 111610 19802
rect 111720 19774 111794 19802
rect 111904 19910 111978 19938
rect 111352 17406 111380 19774
rect 111536 18306 111564 19774
rect 111616 18964 111668 18970
rect 111616 18906 111668 18912
rect 111444 18278 111564 18306
rect 111340 17400 111392 17406
rect 111340 17342 111392 17348
rect 111248 16788 111300 16794
rect 111248 16730 111300 16736
rect 111154 15056 111210 15065
rect 111154 14991 111210 15000
rect 111444 14793 111472 18278
rect 111522 18184 111578 18193
rect 111522 18119 111578 18128
rect 111536 17270 111564 18119
rect 111628 18057 111656 18906
rect 111614 18048 111670 18057
rect 111614 17983 111670 17992
rect 111614 17368 111670 17377
rect 111614 17303 111670 17312
rect 111524 17264 111576 17270
rect 111524 17206 111576 17212
rect 111430 14784 111486 14793
rect 111430 14719 111486 14728
rect 111154 12336 111210 12345
rect 111154 12271 111210 12280
rect 111168 6866 111196 12271
rect 111628 11121 111656 17303
rect 111614 11112 111670 11121
rect 111614 11047 111670 11056
rect 111524 9580 111576 9586
rect 111524 9522 111576 9528
rect 111536 6866 111564 9522
rect 111156 6860 111208 6866
rect 111156 6802 111208 6808
rect 111524 6860 111576 6866
rect 111524 6802 111576 6808
rect 111064 3596 111116 3602
rect 111064 3538 111116 3544
rect 109316 3470 109368 3476
rect 110694 3496 110750 3505
rect 109038 3360 109094 3369
rect 109038 3295 109094 3304
rect 108580 3052 108632 3058
rect 108580 2994 108632 3000
rect 109052 2689 109080 3295
rect 109038 2680 109094 2689
rect 109038 2615 109094 2624
rect 109328 480 109356 3470
rect 110512 3460 110564 3466
rect 110694 3431 110750 3440
rect 110512 3402 110564 3408
rect 110418 2272 110474 2281
rect 110418 2207 110474 2216
rect 110432 814 110460 2207
rect 110420 808 110472 814
rect 110420 750 110472 756
rect 110524 480 110552 3402
rect 111720 3369 111748 19774
rect 111904 17882 111932 19910
rect 111984 19848 112036 19854
rect 112134 19802 112162 20060
rect 111984 19790 112036 19796
rect 111892 17876 111944 17882
rect 111892 17818 111944 17824
rect 111892 15972 111944 15978
rect 111892 15914 111944 15920
rect 111800 11212 111852 11218
rect 111800 11154 111852 11160
rect 111812 9654 111840 11154
rect 111800 9648 111852 9654
rect 111800 9590 111852 9596
rect 111904 6914 111932 15914
rect 111996 9489 112024 19790
rect 112088 19774 112162 19802
rect 112318 19802 112346 20060
rect 112502 19802 112530 20060
rect 112686 19854 112714 20060
rect 112674 19848 112726 19854
rect 112318 19774 112392 19802
rect 112502 19774 112576 19802
rect 112674 19790 112726 19796
rect 112870 19802 112898 20060
rect 113054 19802 113082 20060
rect 113238 19802 113266 20060
rect 112870 19774 112944 19802
rect 111982 9480 112038 9489
rect 111982 9415 112038 9424
rect 111904 6886 112024 6914
rect 111800 4888 111852 4894
rect 111800 4830 111852 4836
rect 111706 3360 111762 3369
rect 111616 3324 111668 3330
rect 111812 3330 111840 4830
rect 111706 3295 111762 3304
rect 111800 3324 111852 3330
rect 111616 3266 111668 3272
rect 111800 3266 111852 3272
rect 111628 480 111656 3266
rect 111798 3224 111854 3233
rect 111798 3159 111854 3168
rect 111812 1329 111840 3159
rect 111798 1320 111854 1329
rect 111798 1255 111854 1264
rect 111996 490 112024 6886
rect 112088 2378 112116 19774
rect 112364 17338 112392 19774
rect 112548 19446 112576 19774
rect 112536 19440 112588 19446
rect 112536 19382 112588 19388
rect 112444 18148 112496 18154
rect 112444 18090 112496 18096
rect 112352 17332 112404 17338
rect 112352 17274 112404 17280
rect 112168 9580 112220 9586
rect 112168 9522 112220 9528
rect 112180 2786 112208 9522
rect 112456 2786 112484 18090
rect 112916 16318 112944 19774
rect 113008 19774 113082 19802
rect 113192 19774 113266 19802
rect 113422 19802 113450 20060
rect 113606 19802 113634 20060
rect 113790 19802 113818 20060
rect 113974 19802 114002 20060
rect 114158 19802 114186 20060
rect 113422 19774 113496 19802
rect 113008 16998 113036 19774
rect 113086 18864 113142 18873
rect 113086 18799 113142 18808
rect 113100 17746 113128 18799
rect 113088 17740 113140 17746
rect 113088 17682 113140 17688
rect 112996 16992 113048 16998
rect 112996 16934 113048 16940
rect 112904 16312 112956 16318
rect 112904 16254 112956 16260
rect 112536 15700 112588 15706
rect 112536 15642 112588 15648
rect 112168 2780 112220 2786
rect 112168 2722 112220 2728
rect 112444 2780 112496 2786
rect 112444 2722 112496 2728
rect 112076 2372 112128 2378
rect 112076 2314 112128 2320
rect 112548 2038 112576 15642
rect 112626 11384 112682 11393
rect 112626 11319 112682 11328
rect 112640 2825 112668 11319
rect 113088 10056 113140 10062
rect 113088 9998 113140 10004
rect 113100 8650 113128 9998
rect 113192 9081 113220 19774
rect 113364 17604 113416 17610
rect 113364 17546 113416 17552
rect 113376 17406 113404 17546
rect 113364 17400 113416 17406
rect 113364 17342 113416 17348
rect 113468 16930 113496 19774
rect 113560 19774 113634 19802
rect 113744 19774 113818 19802
rect 113928 19774 114002 19802
rect 114112 19774 114186 19802
rect 114342 19802 114370 20060
rect 114526 19802 114554 20060
rect 114710 19938 114738 20060
rect 114894 19938 114922 20060
rect 115078 19938 115106 20060
rect 114710 19910 114784 19938
rect 114894 19910 114968 19938
rect 115078 19910 115152 19938
rect 114342 19774 114416 19802
rect 113560 16969 113588 19774
rect 113638 18456 113694 18465
rect 113638 18391 113694 18400
rect 113546 16960 113602 16969
rect 113456 16924 113508 16930
rect 113546 16895 113602 16904
rect 113456 16866 113508 16872
rect 113652 14074 113680 18391
rect 113744 17898 113772 19774
rect 113824 18284 113876 18290
rect 113824 18226 113876 18232
rect 113836 18018 113864 18226
rect 113824 18012 113876 18018
rect 113824 17954 113876 17960
rect 113744 17870 113864 17898
rect 113732 17740 113784 17746
rect 113732 17682 113784 17688
rect 113744 17474 113772 17682
rect 113732 17468 113784 17474
rect 113732 17410 113784 17416
rect 113836 14521 113864 17870
rect 113822 14512 113878 14521
rect 113822 14447 113878 14456
rect 113640 14068 113692 14074
rect 113640 14010 113692 14016
rect 113362 9616 113418 9625
rect 113362 9551 113418 9560
rect 113178 9072 113234 9081
rect 113178 9007 113234 9016
rect 113100 8622 113312 8650
rect 113178 8392 113234 8401
rect 113178 8327 113234 8336
rect 113192 5953 113220 8327
rect 113178 5944 113234 5953
rect 113178 5879 113234 5888
rect 113284 5506 113312 8622
rect 113272 5500 113324 5506
rect 113272 5442 113324 5448
rect 112626 2816 112682 2825
rect 112626 2751 112682 2760
rect 113376 2281 113404 9551
rect 113928 3466 113956 19774
rect 114008 17604 114060 17610
rect 114008 17546 114060 17552
rect 114020 17134 114048 17546
rect 114008 17128 114060 17134
rect 114008 17070 114060 17076
rect 114112 11529 114140 19774
rect 114190 17504 114246 17513
rect 114190 17439 114246 17448
rect 114204 12889 114232 17439
rect 114388 15978 114416 19774
rect 114480 19774 114554 19802
rect 114652 19848 114704 19854
rect 114652 19790 114704 19796
rect 114480 16998 114508 19774
rect 114560 17196 114612 17202
rect 114560 17138 114612 17144
rect 114468 16992 114520 16998
rect 114468 16934 114520 16940
rect 114376 15972 114428 15978
rect 114376 15914 114428 15920
rect 114572 13802 114600 17138
rect 114560 13796 114612 13802
rect 114560 13738 114612 13744
rect 114374 13696 114430 13705
rect 114374 13631 114430 13640
rect 114190 12880 114246 12889
rect 114190 12815 114246 12824
rect 114098 11520 114154 11529
rect 114098 11455 114154 11464
rect 114100 11008 114152 11014
rect 114100 10950 114152 10956
rect 114112 4826 114140 10950
rect 114388 9353 114416 13631
rect 114466 13560 114522 13569
rect 114466 13495 114522 13504
rect 114480 12345 114508 13495
rect 114466 12336 114522 12345
rect 114466 12271 114522 12280
rect 114560 10328 114612 10334
rect 114560 10270 114612 10276
rect 114374 9344 114430 9353
rect 114374 9279 114430 9288
rect 114466 7304 114522 7313
rect 114572 7290 114600 10270
rect 114664 9586 114692 19790
rect 114756 17921 114784 19910
rect 114742 17912 114798 17921
rect 114742 17847 114798 17856
rect 114940 17241 114968 19910
rect 114926 17232 114982 17241
rect 114926 17167 114982 17176
rect 115124 16862 115152 19910
rect 115262 19802 115290 20060
rect 115446 19854 115474 20060
rect 115216 19774 115290 19802
rect 115434 19848 115486 19854
rect 115630 19802 115658 20060
rect 115814 19802 115842 20060
rect 115434 19790 115486 19796
rect 115584 19774 115658 19802
rect 115768 19774 115842 19802
rect 115998 19802 116026 20060
rect 116182 19938 116210 20060
rect 116136 19910 116210 19938
rect 115998 19774 116072 19802
rect 115112 16856 115164 16862
rect 115112 16798 115164 16804
rect 114742 15328 114798 15337
rect 114742 15263 114798 15272
rect 114756 13569 114784 15263
rect 114742 13560 114798 13569
rect 114742 13495 114798 13504
rect 115216 12434 115244 19774
rect 115296 19236 115348 19242
rect 115296 19178 115348 19184
rect 114848 12406 115244 12434
rect 114652 9580 114704 9586
rect 114652 9522 114704 9528
rect 114652 8356 114704 8362
rect 114652 8298 114704 8304
rect 114664 8265 114692 8298
rect 114650 8256 114706 8265
rect 114650 8191 114706 8200
rect 114848 7721 114876 12406
rect 114834 7712 114890 7721
rect 114834 7647 114890 7656
rect 114522 7262 114600 7290
rect 114466 7239 114522 7248
rect 115308 6905 115336 19178
rect 115584 7857 115612 19774
rect 115768 16425 115796 19774
rect 116044 18154 116072 19774
rect 116032 18148 116084 18154
rect 116032 18090 116084 18096
rect 116136 16658 116164 19910
rect 116366 19802 116394 20060
rect 116550 19938 116578 20060
rect 116734 19938 116762 20060
rect 116550 19910 116624 19938
rect 116734 19910 116808 19938
rect 116228 19774 116394 19802
rect 116124 16652 116176 16658
rect 116124 16594 116176 16600
rect 115754 16416 115810 16425
rect 115754 16351 115810 16360
rect 116122 14104 116178 14113
rect 116122 14039 116178 14048
rect 115940 13932 115992 13938
rect 115940 13874 115992 13880
rect 115952 13784 115980 13874
rect 115768 13756 115980 13784
rect 115768 11393 115796 13756
rect 115848 12912 115900 12918
rect 115848 12854 115900 12860
rect 115860 12594 115888 12854
rect 115860 12566 116072 12594
rect 115938 12472 115994 12481
rect 115938 12407 115994 12416
rect 115754 11384 115810 11393
rect 115754 11319 115810 11328
rect 115952 11098 115980 12407
rect 115860 11070 115980 11098
rect 115860 11014 115888 11070
rect 115848 11008 115900 11014
rect 115754 10976 115810 10985
rect 115848 10950 115900 10956
rect 115754 10911 115810 10920
rect 115768 8294 115796 10911
rect 115848 9648 115900 9654
rect 115848 9590 115900 9596
rect 115756 8288 115808 8294
rect 115756 8230 115808 8236
rect 115570 7848 115626 7857
rect 115570 7783 115626 7792
rect 115860 7585 115888 9590
rect 116044 8226 116072 12566
rect 116136 10334 116164 14039
rect 116124 10328 116176 10334
rect 116124 10270 116176 10276
rect 116032 8220 116084 8226
rect 116032 8162 116084 8168
rect 116228 8106 116256 19774
rect 116596 17882 116624 19910
rect 116676 18352 116728 18358
rect 116676 18294 116728 18300
rect 116584 17876 116636 17882
rect 116584 17818 116636 17824
rect 116400 16584 116452 16590
rect 116400 16526 116452 16532
rect 116044 8078 116256 8106
rect 115846 7576 115902 7585
rect 115846 7511 115902 7520
rect 115294 6896 115350 6905
rect 116044 6866 116072 8078
rect 115294 6831 115350 6840
rect 116032 6860 116084 6866
rect 116032 6802 116084 6808
rect 114466 6080 114522 6089
rect 114466 6015 114522 6024
rect 114480 4894 114508 6015
rect 116412 5506 116440 16526
rect 116688 12434 116716 18294
rect 116780 15910 116808 19910
rect 116918 19802 116946 20060
rect 117102 19938 117130 20060
rect 116872 19774 116946 19802
rect 117056 19910 117130 19938
rect 116872 16590 116900 19774
rect 116860 16584 116912 16590
rect 116860 16526 116912 16532
rect 116768 15904 116820 15910
rect 116768 15846 116820 15852
rect 117056 13841 117084 19910
rect 117286 19802 117314 20060
rect 117470 19802 117498 20060
rect 117148 19774 117314 19802
rect 117424 19774 117498 19802
rect 117654 19802 117682 20060
rect 117838 19802 117866 20060
rect 118022 19802 118050 20060
rect 117654 19774 117728 19802
rect 117838 19774 117912 19802
rect 117042 13832 117098 13841
rect 117042 13767 117098 13776
rect 116596 12406 116716 12434
rect 116768 12436 116820 12442
rect 116400 5500 116452 5506
rect 116400 5442 116452 5448
rect 114468 4888 114520 4894
rect 114468 4830 114520 4836
rect 114100 4820 114152 4826
rect 114100 4762 114152 4768
rect 114098 3904 114154 3913
rect 114098 3839 114154 3848
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 113916 3460 113968 3466
rect 113916 3402 113968 3408
rect 113362 2272 113418 2281
rect 113362 2207 113418 2216
rect 112536 2032 112588 2038
rect 112536 1974 112588 1980
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 111996 462 112392 490
rect 114020 480 114048 3538
rect 114112 1222 114140 3839
rect 115204 3664 115256 3670
rect 115204 3606 115256 3612
rect 114468 2780 114520 2786
rect 114468 2722 114520 2728
rect 114480 1290 114508 2722
rect 114468 1284 114520 1290
rect 114468 1226 114520 1232
rect 114100 1216 114152 1222
rect 114100 1158 114152 1164
rect 115216 480 115244 3606
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 115848 2848 115900 2854
rect 115848 2790 115900 2796
rect 115860 2689 115888 2790
rect 115846 2680 115902 2689
rect 115846 2615 115902 2624
rect 115848 1896 115900 1902
rect 115848 1838 115900 1844
rect 115860 1358 115888 1838
rect 115848 1352 115900 1358
rect 115848 1294 115900 1300
rect 116412 480 116440 3470
rect 116596 2650 116624 12406
rect 116768 12378 116820 12384
rect 116780 11150 116808 12378
rect 116768 11144 116820 11150
rect 116768 11086 116820 11092
rect 117148 9353 117176 19774
rect 117424 19718 117452 19774
rect 117412 19712 117464 19718
rect 117412 19654 117464 19660
rect 117410 17912 117466 17921
rect 117410 17847 117466 17856
rect 117320 16516 117372 16522
rect 117320 16458 117372 16464
rect 117332 16318 117360 16458
rect 117228 16312 117280 16318
rect 117228 16254 117280 16260
rect 117320 16312 117372 16318
rect 117320 16254 117372 16260
rect 117240 13569 117268 16254
rect 117424 15337 117452 17847
rect 117700 17474 117728 19774
rect 117884 17882 117912 19774
rect 117976 19774 118050 19802
rect 118206 19802 118234 20060
rect 118390 19802 118418 20060
rect 118574 19802 118602 20060
rect 118206 19774 118280 19802
rect 117872 17876 117924 17882
rect 117872 17818 117924 17824
rect 117688 17468 117740 17474
rect 117688 17410 117740 17416
rect 117688 17060 117740 17066
rect 117688 17002 117740 17008
rect 117504 16856 117556 16862
rect 117504 16798 117556 16804
rect 117410 15328 117466 15337
rect 117410 15263 117466 15272
rect 117226 13560 117282 13569
rect 117226 13495 117282 13504
rect 117516 13025 117544 16798
rect 117594 15464 117650 15473
rect 117594 15399 117650 15408
rect 117502 13016 117558 13025
rect 117502 12951 117558 12960
rect 117608 10849 117636 15399
rect 117700 14074 117728 17002
rect 117688 14068 117740 14074
rect 117688 14010 117740 14016
rect 117976 13938 118004 19774
rect 118054 18048 118110 18057
rect 118054 17983 118110 17992
rect 117964 13932 118016 13938
rect 117964 13874 118016 13880
rect 118068 13818 118096 17983
rect 118252 17950 118280 19774
rect 118344 19774 118418 19802
rect 118528 19774 118602 19802
rect 118758 19802 118786 20060
rect 118942 19802 118970 20060
rect 119126 19802 119154 20060
rect 119310 19802 119338 20060
rect 118758 19774 118832 19802
rect 118942 19774 119016 19802
rect 118240 17944 118292 17950
rect 118240 17886 118292 17892
rect 118148 15768 118200 15774
rect 118148 15710 118200 15716
rect 117976 13790 118096 13818
rect 117594 10840 117650 10849
rect 117594 10775 117650 10784
rect 117134 9344 117190 9353
rect 117134 9279 117190 9288
rect 116676 4140 116728 4146
rect 116676 4082 116728 4088
rect 116688 3670 116716 4082
rect 116676 3664 116728 3670
rect 116676 3606 116728 3612
rect 117872 3596 117924 3602
rect 117872 3538 117924 3544
rect 117884 3330 117912 3538
rect 117872 3324 117924 3330
rect 117872 3266 117924 3272
rect 117596 3188 117648 3194
rect 117596 3130 117648 3136
rect 116584 2644 116636 2650
rect 116584 2586 116636 2592
rect 117608 480 117636 3130
rect 117872 2644 117924 2650
rect 117872 2586 117924 2592
rect 112364 354 112392 462
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 117884 474 117912 2586
rect 117976 2553 118004 13790
rect 118056 12912 118108 12918
rect 118056 12854 118108 12860
rect 118068 4894 118096 12854
rect 118056 4888 118108 4894
rect 118056 4830 118108 4836
rect 118160 2553 118188 15710
rect 118344 13705 118372 19774
rect 118424 19372 118476 19378
rect 118424 19314 118476 19320
rect 118330 13696 118386 13705
rect 118330 13631 118386 13640
rect 118238 13560 118294 13569
rect 118238 13495 118294 13504
rect 118252 3534 118280 13495
rect 118436 12918 118464 19314
rect 118528 18601 118556 19774
rect 118514 18592 118570 18601
rect 118514 18527 118570 18536
rect 118698 17776 118754 17785
rect 118804 17762 118832 19774
rect 118804 17734 118924 17762
rect 118698 17711 118754 17720
rect 118712 13818 118740 17711
rect 118790 17640 118846 17649
rect 118790 17575 118846 17584
rect 118804 14113 118832 17575
rect 118896 17270 118924 17734
rect 118884 17264 118936 17270
rect 118884 17206 118936 17212
rect 118988 15065 119016 19774
rect 119080 19774 119154 19802
rect 119264 19774 119338 19802
rect 119494 19802 119522 20060
rect 119678 19802 119706 20060
rect 119862 19922 119890 20060
rect 119850 19916 119902 19922
rect 119850 19858 119902 19864
rect 120046 19802 120074 20060
rect 120230 19802 120258 20060
rect 119494 19774 119568 19802
rect 119080 17513 119108 19774
rect 119066 17504 119122 17513
rect 119066 17439 119122 17448
rect 118974 15056 119030 15065
rect 118974 14991 119030 15000
rect 118790 14104 118846 14113
rect 118790 14039 118846 14048
rect 118792 13932 118844 13938
rect 118792 13874 118844 13880
rect 118620 13790 118740 13818
rect 118804 13802 118832 13874
rect 118792 13796 118844 13802
rect 118424 12912 118476 12918
rect 118424 12854 118476 12860
rect 118620 12481 118648 13790
rect 118792 13738 118844 13744
rect 118606 12472 118662 12481
rect 118606 12407 118662 12416
rect 119264 10985 119292 19774
rect 119344 19168 119396 19174
rect 119344 19110 119396 19116
rect 119250 10976 119306 10985
rect 119250 10911 119306 10920
rect 119356 8294 119384 19110
rect 119540 17762 119568 19774
rect 119632 19774 119706 19802
rect 120000 19774 120074 19802
rect 120184 19774 120258 19802
rect 120414 19802 120442 20060
rect 120598 19802 120626 20060
rect 120782 19802 120810 20060
rect 120414 19774 120488 19802
rect 119632 17921 119660 19774
rect 119618 17912 119674 17921
rect 119618 17847 119674 17856
rect 119802 17912 119858 17921
rect 119802 17847 119858 17856
rect 119816 17762 119844 17847
rect 119540 17734 119844 17762
rect 119528 17468 119580 17474
rect 119528 17410 119580 17416
rect 119540 12986 119568 17410
rect 119896 14068 119948 14074
rect 119896 14010 119948 14016
rect 119436 12980 119488 12986
rect 119436 12922 119488 12928
rect 119528 12980 119580 12986
rect 119528 12922 119580 12928
rect 119344 8288 119396 8294
rect 119344 8230 119396 8236
rect 118698 6896 118754 6905
rect 118698 6831 118700 6840
rect 118752 6831 118754 6840
rect 118700 6802 118752 6808
rect 119448 4146 119476 12922
rect 119908 9761 119936 14010
rect 120000 12209 120028 19774
rect 120080 18352 120132 18358
rect 120080 18294 120132 18300
rect 119986 12200 120042 12209
rect 119986 12135 120042 12144
rect 119894 9752 119950 9761
rect 119894 9687 119950 9696
rect 120092 9625 120120 18294
rect 120184 17785 120212 19774
rect 120170 17776 120226 17785
rect 120170 17711 120226 17720
rect 120460 17474 120488 19774
rect 120552 19774 120626 19802
rect 120736 19774 120810 19802
rect 120966 19802 120994 20060
rect 121150 19802 121178 20060
rect 121334 19825 121362 20060
rect 120966 19774 121040 19802
rect 120448 17468 120500 17474
rect 120448 17410 120500 17416
rect 120078 9616 120134 9625
rect 120078 9551 120134 9560
rect 119896 8220 119948 8226
rect 119896 8162 119948 8168
rect 119436 4140 119488 4146
rect 119436 4082 119488 4088
rect 118240 3528 118292 3534
rect 118240 3470 118292 3476
rect 118792 3256 118844 3262
rect 118792 3198 118844 3204
rect 118608 2916 118660 2922
rect 118608 2858 118660 2864
rect 117962 2544 118018 2553
rect 117962 2479 118018 2488
rect 118146 2544 118202 2553
rect 118620 2514 118648 2858
rect 118146 2479 118202 2488
rect 118608 2508 118660 2514
rect 118608 2450 118660 2456
rect 118804 480 118832 3198
rect 119908 480 119936 8162
rect 120552 7721 120580 19774
rect 120736 18358 120764 19774
rect 121012 19281 121040 19774
rect 121104 19774 121178 19802
rect 121320 19816 121376 19825
rect 120998 19272 121054 19281
rect 120998 19207 121054 19216
rect 120724 18352 120776 18358
rect 120724 18294 120776 18300
rect 121000 18284 121052 18290
rect 121000 18226 121052 18232
rect 120724 18012 120776 18018
rect 120724 17954 120776 17960
rect 120538 7712 120594 7721
rect 120538 7647 120594 7656
rect 120736 2378 120764 17954
rect 120908 17264 120960 17270
rect 120908 17206 120960 17212
rect 120920 16930 120948 17206
rect 120908 16924 120960 16930
rect 120908 16866 120960 16872
rect 120814 16688 120870 16697
rect 120814 16623 120870 16632
rect 120828 5953 120856 16623
rect 121012 6866 121040 18226
rect 121104 16017 121132 19774
rect 121518 19802 121546 20060
rect 121702 19802 121730 20060
rect 121886 19802 121914 20060
rect 121320 19751 121376 19760
rect 121472 19774 121546 19802
rect 121656 19774 121730 19802
rect 121840 19774 121914 19802
rect 122070 19802 122098 20060
rect 122254 19802 122282 20060
rect 122438 19802 122466 20060
rect 122070 19774 122144 19802
rect 121368 17944 121420 17950
rect 121368 17886 121420 17892
rect 121276 17876 121328 17882
rect 121276 17818 121328 17824
rect 121184 16584 121236 16590
rect 121184 16526 121236 16532
rect 121090 16008 121146 16017
rect 121090 15943 121146 15952
rect 121000 6860 121052 6866
rect 121000 6802 121052 6808
rect 120814 5944 120870 5953
rect 120814 5879 120870 5888
rect 121196 4894 121224 16526
rect 121288 9489 121316 17818
rect 121380 12753 121408 17886
rect 121366 12744 121422 12753
rect 121366 12679 121422 12688
rect 121274 9480 121330 9489
rect 121274 9415 121330 9424
rect 121276 7472 121328 7478
rect 121276 7414 121328 7420
rect 121184 4888 121236 4894
rect 121184 4830 121236 4836
rect 121288 3398 121316 7414
rect 121472 4826 121500 19774
rect 121552 19644 121604 19650
rect 121552 19586 121604 19592
rect 121564 19106 121592 19586
rect 121552 19100 121604 19106
rect 121552 19042 121604 19048
rect 121552 18012 121604 18018
rect 121552 17954 121604 17960
rect 121564 15473 121592 17954
rect 121550 15464 121606 15473
rect 121550 15399 121606 15408
rect 121656 5001 121684 19774
rect 121840 18057 121868 19774
rect 122116 19689 122144 19774
rect 122208 19774 122282 19802
rect 122392 19774 122466 19802
rect 122622 19802 122650 20060
rect 122806 19802 122834 20060
rect 122990 19802 123018 20060
rect 122622 19774 122696 19802
rect 122102 19680 122158 19689
rect 122012 19644 122064 19650
rect 122102 19615 122158 19624
rect 122012 19586 122064 19592
rect 121920 19372 121972 19378
rect 121920 19314 121972 19320
rect 121932 19174 121960 19314
rect 121920 19168 121972 19174
rect 121920 19110 121972 19116
rect 121826 18048 121882 18057
rect 121826 17983 121882 17992
rect 121736 17128 121788 17134
rect 121736 17070 121788 17076
rect 121748 13938 121776 17070
rect 122024 15201 122052 19586
rect 122104 19372 122156 19378
rect 122104 19314 122156 19320
rect 122010 15192 122066 15201
rect 122010 15127 122066 15136
rect 121736 13932 121788 13938
rect 121736 13874 121788 13880
rect 121642 4992 121698 5001
rect 121642 4927 121698 4936
rect 121460 4820 121512 4826
rect 121460 4762 121512 4768
rect 121092 3392 121144 3398
rect 121092 3334 121144 3340
rect 121276 3392 121328 3398
rect 121276 3334 121328 3340
rect 120724 2372 120776 2378
rect 120724 2314 120776 2320
rect 121104 480 121132 3334
rect 122116 2417 122144 19314
rect 122208 13802 122236 19774
rect 122392 17649 122420 19774
rect 122472 19032 122524 19038
rect 122472 18974 122524 18980
rect 122378 17640 122434 17649
rect 122378 17575 122434 17584
rect 122288 17468 122340 17474
rect 122288 17410 122340 17416
rect 122380 17468 122432 17474
rect 122380 17410 122432 17416
rect 122300 15162 122328 17410
rect 122392 16998 122420 17410
rect 122380 16992 122432 16998
rect 122380 16934 122432 16940
rect 122378 15328 122434 15337
rect 122378 15263 122434 15272
rect 122288 15156 122340 15162
rect 122288 15098 122340 15104
rect 122196 13796 122248 13802
rect 122196 13738 122248 13744
rect 122392 3913 122420 15263
rect 122484 8226 122512 18974
rect 122668 16658 122696 19774
rect 122760 19774 122834 19802
rect 122944 19774 123018 19802
rect 123174 19802 123202 20060
rect 123358 19802 123386 20060
rect 123174 19774 123248 19802
rect 122656 16652 122708 16658
rect 122656 16594 122708 16600
rect 122760 15774 122788 19774
rect 122838 17640 122894 17649
rect 122838 17575 122894 17584
rect 122748 15768 122800 15774
rect 122748 15710 122800 15716
rect 122852 13433 122880 17575
rect 122944 16833 122972 19774
rect 123022 18592 123078 18601
rect 123022 18527 123078 18536
rect 122930 16824 122986 16833
rect 122930 16759 122986 16768
rect 123036 15337 123064 18527
rect 123116 18352 123168 18358
rect 123116 18294 123168 18300
rect 123128 17921 123156 18294
rect 123220 17950 123248 19774
rect 123312 19774 123386 19802
rect 123542 19802 123570 20060
rect 123726 19802 123754 20060
rect 123910 19802 123938 20060
rect 124094 19802 124122 20060
rect 124278 19802 124306 20060
rect 124462 19802 124490 20060
rect 124646 19802 124674 20060
rect 123542 19774 123616 19802
rect 123208 17944 123260 17950
rect 123114 17912 123170 17921
rect 123208 17886 123260 17892
rect 123114 17847 123170 17856
rect 123022 15328 123078 15337
rect 123022 15263 123078 15272
rect 123312 13938 123340 19774
rect 123482 17912 123538 17921
rect 123482 17847 123538 17856
rect 123300 13932 123352 13938
rect 123300 13874 123352 13880
rect 122838 13424 122894 13433
rect 122838 13359 122894 13368
rect 123496 9722 123524 17847
rect 123588 16697 123616 19774
rect 123680 19774 123754 19802
rect 123864 19774 123938 19802
rect 124048 19774 124122 19802
rect 124232 19774 124306 19802
rect 124416 19774 124490 19802
rect 124600 19774 124674 19802
rect 124830 19802 124858 20060
rect 125014 19802 125042 20060
rect 125198 19802 125226 20060
rect 125382 19802 125410 20060
rect 125566 19802 125594 20060
rect 125750 19802 125778 20060
rect 125934 19802 125962 20060
rect 124830 19774 124904 19802
rect 123574 16688 123630 16697
rect 123574 16623 123630 16632
rect 123576 15768 123628 15774
rect 123576 15710 123628 15716
rect 123484 9716 123536 9722
rect 123484 9658 123536 9664
rect 123024 8288 123076 8294
rect 123024 8230 123076 8236
rect 122472 8220 122524 8226
rect 122472 8162 122524 8168
rect 122378 3904 122434 3913
rect 122378 3839 122434 3848
rect 122288 2916 122340 2922
rect 122288 2858 122340 2864
rect 122102 2408 122158 2417
rect 122102 2343 122158 2352
rect 121460 1964 121512 1970
rect 121460 1906 121512 1912
rect 121184 1692 121236 1698
rect 121184 1634 121236 1640
rect 121196 1358 121224 1634
rect 121368 1624 121420 1630
rect 121368 1566 121420 1572
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 121380 1290 121408 1566
rect 121472 1290 121500 1906
rect 121368 1284 121420 1290
rect 121368 1226 121420 1232
rect 121460 1284 121512 1290
rect 121460 1226 121512 1232
rect 122300 480 122328 2858
rect 122840 1556 122892 1562
rect 122840 1498 122892 1504
rect 122748 1488 122800 1494
rect 122748 1430 122800 1436
rect 122760 950 122788 1430
rect 122852 1329 122880 1498
rect 123036 1426 123064 8230
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 122932 1420 122984 1426
rect 122932 1362 122984 1368
rect 123024 1420 123076 1426
rect 123024 1362 123076 1368
rect 122838 1320 122894 1329
rect 122838 1255 122894 1264
rect 122944 950 122972 1362
rect 122748 944 122800 950
rect 122748 886 122800 892
rect 122932 944 122984 950
rect 122932 886 122984 892
rect 123496 480 123524 4082
rect 123588 2417 123616 15710
rect 123680 13841 123708 19774
rect 123760 16652 123812 16658
rect 123760 16594 123812 16600
rect 123666 13832 123722 13841
rect 123666 13767 123722 13776
rect 123772 9654 123800 16594
rect 123864 16574 123892 19774
rect 124048 18018 124076 19774
rect 124036 18012 124088 18018
rect 124036 17954 124088 17960
rect 124232 17921 124260 19774
rect 124312 18148 124364 18154
rect 124312 18090 124364 18096
rect 124218 17912 124274 17921
rect 124218 17847 124274 17856
rect 123864 16546 124260 16574
rect 124128 15156 124180 15162
rect 124128 15098 124180 15104
rect 124140 11121 124168 15098
rect 124232 13977 124260 16546
rect 124324 15230 124352 18090
rect 124312 15224 124364 15230
rect 124416 15201 124444 19774
rect 124600 19174 124628 19774
rect 124588 19168 124640 19174
rect 124588 19110 124640 19116
rect 124876 19038 124904 19774
rect 124968 19774 125042 19802
rect 125152 19774 125226 19802
rect 125336 19774 125410 19802
rect 125520 19774 125594 19802
rect 125704 19774 125778 19802
rect 125888 19774 125962 19802
rect 126118 19802 126146 20060
rect 126302 19802 126330 20060
rect 126486 19802 126514 20060
rect 126118 19774 126192 19802
rect 124968 19378 124996 19774
rect 124956 19372 125008 19378
rect 124956 19314 125008 19320
rect 124864 19032 124916 19038
rect 124864 18974 124916 18980
rect 125152 18465 125180 19774
rect 125138 18456 125194 18465
rect 125138 18391 125194 18400
rect 125046 17912 125102 17921
rect 125046 17847 125102 17856
rect 124862 17776 124918 17785
rect 124862 17711 124918 17720
rect 124312 15166 124364 15172
rect 124402 15192 124458 15201
rect 124402 15127 124458 15136
rect 124218 13968 124274 13977
rect 124218 13903 124274 13912
rect 124218 13832 124274 13841
rect 124218 13767 124274 13776
rect 124126 11112 124182 11121
rect 124126 11047 124182 11056
rect 123760 9648 123812 9654
rect 123760 9590 123812 9596
rect 124232 8945 124260 13767
rect 124588 9648 124640 9654
rect 124588 9590 124640 9596
rect 124218 8936 124274 8945
rect 124218 8871 124274 8880
rect 124220 7540 124272 7546
rect 124220 7482 124272 7488
rect 124232 2650 124260 7482
rect 124600 3194 124628 9590
rect 124680 4072 124732 4078
rect 124680 4014 124732 4020
rect 124588 3188 124640 3194
rect 124588 3130 124640 3136
rect 124220 2644 124272 2650
rect 124220 2586 124272 2592
rect 123574 2408 123630 2417
rect 123574 2343 123630 2352
rect 124128 1692 124180 1698
rect 124128 1634 124180 1640
rect 124140 1601 124168 1634
rect 124126 1592 124182 1601
rect 124126 1527 124182 1536
rect 123680 882 123892 898
rect 123668 876 123904 882
rect 123720 870 123852 876
rect 123668 818 123720 824
rect 123852 818 123904 824
rect 124692 480 124720 4014
rect 124876 1562 124904 17711
rect 125060 8362 125088 17847
rect 125336 13433 125364 19774
rect 125520 17513 125548 19774
rect 125704 17921 125732 19774
rect 125690 17912 125746 17921
rect 125690 17847 125746 17856
rect 125506 17504 125562 17513
rect 125506 17439 125562 17448
rect 125508 13864 125560 13870
rect 125888 13841 125916 19774
rect 126164 17066 126192 19774
rect 126256 19774 126330 19802
rect 126440 19774 126514 19802
rect 126670 19802 126698 20060
rect 126854 19802 126882 20060
rect 126670 19774 126744 19802
rect 126256 17785 126284 19774
rect 126242 17776 126298 17785
rect 126242 17711 126298 17720
rect 126152 17060 126204 17066
rect 126152 17002 126204 17008
rect 126242 15056 126298 15065
rect 126242 14991 126298 15000
rect 125508 13806 125560 13812
rect 125874 13832 125930 13841
rect 125322 13424 125378 13433
rect 125322 13359 125378 13368
rect 125520 12322 125548 13806
rect 125874 13767 125930 13776
rect 125520 12294 125640 12322
rect 125140 11552 125192 11558
rect 125140 11494 125192 11500
rect 125152 9858 125180 11494
rect 125140 9852 125192 9858
rect 125140 9794 125192 9800
rect 125048 8356 125100 8362
rect 125048 8298 125100 8304
rect 125612 7886 125640 12294
rect 126256 12073 126284 14991
rect 126242 12064 126298 12073
rect 126242 11999 126298 12008
rect 125600 7880 125652 7886
rect 125600 7822 125652 7828
rect 124864 1556 124916 1562
rect 124864 1498 124916 1504
rect 125876 1488 125928 1494
rect 125876 1430 125928 1436
rect 125888 480 125916 1430
rect 117872 468 117924 474
rect 117872 410 117924 416
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126440 105 126468 19774
rect 126716 19689 126744 19774
rect 126808 19774 126882 19802
rect 127038 19802 127066 20060
rect 127222 19802 127250 20060
rect 127406 19938 127434 20060
rect 127360 19910 127434 19938
rect 127038 19774 127112 19802
rect 127222 19774 127296 19802
rect 126702 19680 126758 19689
rect 126808 19650 126836 19774
rect 126702 19615 126758 19624
rect 126796 19644 126848 19650
rect 126796 19586 126848 19592
rect 126520 17944 126572 17950
rect 126520 17886 126572 17892
rect 126532 13870 126560 17886
rect 126888 17196 126940 17202
rect 126888 17138 126940 17144
rect 126900 16561 126928 17138
rect 126886 16552 126942 16561
rect 126886 16487 126942 16496
rect 126520 13864 126572 13870
rect 126520 13806 126572 13812
rect 126886 11520 126942 11529
rect 126886 11455 126942 11464
rect 126900 10985 126928 11455
rect 126886 10976 126942 10985
rect 126886 10911 126942 10920
rect 127084 2689 127112 19774
rect 127268 19553 127296 19774
rect 127254 19544 127310 19553
rect 127254 19479 127310 19488
rect 127360 17649 127388 19910
rect 127440 19848 127492 19854
rect 127440 19790 127492 19796
rect 127590 19802 127618 20060
rect 127774 19802 127802 20060
rect 127958 19938 127986 20060
rect 127958 19910 128032 19938
rect 127452 19378 127480 19790
rect 127590 19774 127664 19802
rect 127440 19372 127492 19378
rect 127440 19314 127492 19320
rect 127636 17921 127664 19774
rect 127728 19774 127802 19802
rect 127900 19848 127952 19854
rect 127900 19790 127952 19796
rect 127622 17912 127678 17921
rect 127622 17847 127678 17856
rect 127346 17640 127402 17649
rect 127346 17575 127402 17584
rect 127624 13864 127676 13870
rect 127624 13806 127676 13812
rect 127532 9852 127584 9858
rect 127532 9794 127584 9800
rect 127544 6934 127572 9794
rect 127532 6928 127584 6934
rect 127532 6870 127584 6876
rect 127636 5982 127664 13806
rect 127728 7585 127756 19774
rect 127912 19281 127940 19790
rect 127898 19272 127954 19281
rect 127898 19207 127954 19216
rect 128004 18601 128032 19910
rect 128142 19802 128170 20060
rect 128326 19802 128354 20060
rect 128142 19774 128216 19802
rect 128188 19174 128216 19774
rect 128280 19774 128354 19802
rect 128510 19802 128538 20060
rect 128694 19802 128722 20060
rect 128878 19802 128906 20060
rect 128510 19774 128584 19802
rect 128694 19774 128768 19802
rect 128176 19168 128228 19174
rect 128176 19110 128228 19116
rect 127990 18592 128046 18601
rect 127990 18527 128046 18536
rect 128280 16833 128308 19774
rect 128452 19644 128504 19650
rect 128452 19586 128504 19592
rect 128360 19032 128412 19038
rect 128360 18974 128412 18980
rect 128372 18601 128400 18974
rect 128358 18592 128414 18601
rect 128358 18527 128414 18536
rect 128464 18358 128492 19586
rect 128556 19038 128584 19774
rect 128544 19032 128596 19038
rect 128544 18974 128596 18980
rect 128452 18352 128504 18358
rect 128452 18294 128504 18300
rect 128360 18284 128412 18290
rect 128360 18226 128412 18232
rect 128266 16824 128322 16833
rect 128266 16759 128322 16768
rect 127808 7880 127860 7886
rect 127808 7822 127860 7828
rect 127714 7576 127770 7585
rect 127714 7511 127770 7520
rect 127624 5976 127676 5982
rect 127624 5918 127676 5924
rect 127624 4616 127676 4622
rect 127624 4558 127676 4564
rect 127636 4146 127664 4558
rect 127624 4140 127676 4146
rect 127624 4082 127676 4088
rect 127820 4078 127848 7822
rect 128372 6914 128400 18226
rect 128740 17785 128768 19774
rect 128832 19774 128906 19802
rect 129062 19802 129090 20060
rect 129246 19802 129274 20060
rect 129430 19802 129458 20060
rect 129614 19802 129642 20060
rect 129798 19802 129826 20060
rect 129982 19802 130010 20060
rect 129062 19774 129136 19802
rect 129246 19774 129320 19802
rect 129430 19774 129504 19802
rect 129614 19774 129688 19802
rect 129798 19774 129872 19802
rect 128726 17776 128782 17785
rect 128726 17711 128782 17720
rect 128832 16425 128860 19774
rect 129108 18562 129136 19774
rect 129096 18556 129148 18562
rect 129096 18498 129148 18504
rect 129292 17921 129320 19774
rect 128910 17912 128966 17921
rect 128910 17847 128966 17856
rect 129278 17912 129334 17921
rect 129278 17847 129334 17856
rect 128818 16416 128874 16425
rect 128818 16351 128874 16360
rect 128544 15224 128596 15230
rect 128544 15166 128596 15172
rect 128452 10260 128504 10266
rect 128452 10202 128504 10208
rect 128464 8702 128492 10202
rect 128556 10062 128584 15166
rect 128924 10849 128952 17847
rect 129476 17649 129504 19774
rect 129556 19100 129608 19106
rect 129556 19042 129608 19048
rect 129462 17640 129518 17649
rect 129462 17575 129518 17584
rect 129568 16590 129596 19042
rect 129660 19009 129688 19774
rect 129646 19000 129702 19009
rect 129646 18935 129702 18944
rect 129740 16652 129792 16658
rect 129740 16594 129792 16600
rect 129556 16584 129608 16590
rect 129752 16561 129780 16594
rect 129556 16526 129608 16532
rect 129738 16552 129794 16561
rect 129738 16487 129794 16496
rect 129844 15745 129872 19774
rect 129936 19774 130010 19802
rect 130166 19802 130194 20060
rect 130350 19802 130378 20060
rect 130534 19802 130562 20060
rect 150624 19848 150676 19854
rect 130166 19774 130240 19802
rect 130350 19774 130424 19802
rect 130534 19774 130608 19802
rect 150624 19790 150676 19796
rect 129830 15736 129886 15745
rect 129830 15671 129886 15680
rect 129740 13932 129792 13938
rect 129740 13874 129792 13880
rect 129002 13832 129058 13841
rect 129002 13767 129058 13776
rect 128910 10840 128966 10849
rect 128910 10775 128966 10784
rect 128544 10056 128596 10062
rect 128544 9998 128596 10004
rect 128452 8696 128504 8702
rect 128452 8638 128504 8644
rect 128372 6886 128952 6914
rect 127808 4072 127860 4078
rect 127808 4014 127860 4020
rect 128176 3392 128228 3398
rect 128176 3334 128228 3340
rect 127070 2680 127126 2689
rect 127070 2615 127126 2624
rect 126978 1592 127034 1601
rect 126978 1527 127034 1536
rect 126992 1358 127020 1527
rect 126980 1352 127032 1358
rect 126980 1294 127032 1300
rect 128188 480 128216 3334
rect 128360 1624 128412 1630
rect 128360 1566 128412 1572
rect 128372 814 128400 1566
rect 128360 808 128412 814
rect 128360 750 128412 756
rect 126426 96 126482 105
rect 126950 82 127062 480
rect 126624 66 127062 82
rect 126426 31 126482 40
rect 126612 60 127062 66
rect 126664 54 127062 60
rect 126612 2 126664 8
rect 126950 -960 127062 54
rect 128146 -960 128258 480
rect 128924 354 128952 6886
rect 129016 4729 129044 13767
rect 129752 7886 129780 13874
rect 129740 7880 129792 7886
rect 129740 7822 129792 7828
rect 129936 4865 129964 19774
rect 130014 17776 130070 17785
rect 130014 17711 130070 17720
rect 130028 15230 130056 17711
rect 130212 17377 130240 19774
rect 130198 17368 130254 17377
rect 130198 17303 130254 17312
rect 130396 17241 130424 19774
rect 130580 17785 130608 19774
rect 149060 19712 149112 19718
rect 149060 19654 149112 19660
rect 142620 19644 142672 19650
rect 142620 19586 142672 19592
rect 131120 19576 131172 19582
rect 131120 19518 131172 19524
rect 131132 19106 131160 19518
rect 142632 19281 142660 19586
rect 148324 19508 148376 19514
rect 148324 19450 148376 19456
rect 142618 19272 142674 19281
rect 142618 19207 142674 19216
rect 131120 19100 131172 19106
rect 131120 19042 131172 19048
rect 147680 19032 147732 19038
rect 137282 19000 137338 19009
rect 147680 18974 147732 18980
rect 137282 18935 137338 18944
rect 135352 18896 135404 18902
rect 135352 18838 135404 18844
rect 130658 17912 130714 17921
rect 130658 17847 130714 17856
rect 130566 17776 130622 17785
rect 130566 17711 130622 17720
rect 130382 17232 130438 17241
rect 130382 17167 130438 17176
rect 130016 15224 130068 15230
rect 130016 15166 130068 15172
rect 130292 8288 130344 8294
rect 130292 8230 130344 8236
rect 129922 4856 129978 4865
rect 129922 4791 129978 4800
rect 129002 4720 129058 4729
rect 129002 4655 129058 4664
rect 129740 2916 129792 2922
rect 129740 2858 129792 2864
rect 129752 2038 129780 2858
rect 129740 2032 129792 2038
rect 129740 1974 129792 1980
rect 129646 1320 129702 1329
rect 129646 1255 129648 1264
rect 129700 1255 129702 1264
rect 129648 1226 129700 1232
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130304 66 130332 8230
rect 130672 5681 130700 17847
rect 131120 17060 131172 17066
rect 131120 17002 131172 17008
rect 131132 16561 131160 17002
rect 132500 16652 132552 16658
rect 132500 16594 132552 16600
rect 131118 16552 131174 16561
rect 131118 16487 131174 16496
rect 131118 15736 131174 15745
rect 132512 15706 132540 16594
rect 133788 16584 133840 16590
rect 133788 16526 133840 16532
rect 131118 15671 131174 15680
rect 132500 15700 132552 15706
rect 131132 15026 131160 15671
rect 132500 15642 132552 15648
rect 131120 15020 131172 15026
rect 131120 14962 131172 14968
rect 131304 14408 131356 14414
rect 131304 14350 131356 14356
rect 131120 10192 131172 10198
rect 131120 10134 131172 10140
rect 131132 9722 131160 10134
rect 131120 9716 131172 9722
rect 131120 9658 131172 9664
rect 131212 8696 131264 8702
rect 131212 8638 131264 8644
rect 130658 5672 130714 5681
rect 130658 5607 130714 5616
rect 131120 4616 131172 4622
rect 131120 4558 131172 4564
rect 131132 4146 131160 4558
rect 131120 4140 131172 4146
rect 131120 4082 131172 4088
rect 131224 3398 131252 8638
rect 131212 3392 131264 3398
rect 131212 3334 131264 3340
rect 130568 2644 130620 2650
rect 130568 2586 130620 2592
rect 130580 480 130608 2586
rect 130292 60 130344 66
rect 130292 2 130344 8
rect 130538 -960 130650 480
rect 131316 354 131344 14350
rect 132590 13696 132646 13705
rect 132590 13631 132646 13640
rect 132604 10334 132632 13631
rect 133800 12578 133828 16526
rect 133788 12572 133840 12578
rect 133788 12514 133840 12520
rect 133236 11348 133288 11354
rect 133236 11290 133288 11296
rect 133248 10985 133276 11290
rect 133234 10976 133290 10985
rect 133234 10911 133290 10920
rect 132592 10328 132644 10334
rect 132592 10270 132644 10276
rect 135168 10124 135220 10130
rect 135168 10066 135220 10072
rect 135180 8838 135208 10066
rect 135168 8832 135220 8838
rect 135168 8774 135220 8780
rect 134156 6928 134208 6934
rect 135364 6914 135392 18838
rect 136088 18012 136140 18018
rect 136088 17954 136140 17960
rect 136100 11354 136128 17954
rect 137296 17950 137324 18935
rect 146944 18556 146996 18562
rect 146944 18498 146996 18504
rect 143446 18184 143502 18193
rect 143446 18119 143502 18128
rect 137284 17944 137336 17950
rect 137284 17886 137336 17892
rect 143460 17882 143488 18119
rect 146208 18012 146260 18018
rect 146208 17954 146260 17960
rect 143448 17876 143500 17882
rect 143448 17818 143500 17824
rect 146220 17649 146248 17954
rect 142250 17640 142306 17649
rect 142250 17575 142306 17584
rect 146206 17640 146262 17649
rect 146206 17575 146262 17584
rect 142160 17196 142212 17202
rect 142160 17138 142212 17144
rect 142172 16590 142200 17138
rect 142160 16584 142212 16590
rect 142160 16526 142212 16532
rect 142264 15094 142292 17575
rect 143538 17504 143594 17513
rect 143538 17439 143594 17448
rect 143552 16522 143580 17439
rect 143632 17196 143684 17202
rect 143632 17138 143684 17144
rect 143540 16516 143592 16522
rect 143540 16458 143592 16464
rect 143644 15842 143672 17138
rect 146300 17060 146352 17066
rect 146300 17002 146352 17008
rect 146312 16574 146340 17002
rect 146312 16546 146892 16574
rect 143632 15836 143684 15842
rect 143632 15778 143684 15784
rect 143080 15700 143132 15706
rect 143080 15642 143132 15648
rect 142252 15088 142304 15094
rect 142252 15030 142304 15036
rect 137284 13864 137336 13870
rect 137284 13806 137336 13812
rect 137296 13705 137324 13806
rect 137282 13696 137338 13705
rect 137282 13631 137338 13640
rect 140136 12572 140188 12578
rect 140136 12514 140188 12520
rect 136088 11348 136140 11354
rect 136088 11290 136140 11296
rect 139308 8832 139360 8838
rect 139308 8774 139360 8780
rect 137928 8288 137980 8294
rect 137928 8230 137980 8236
rect 135364 6886 136496 6914
rect 134156 6870 134208 6876
rect 133788 4684 133840 4690
rect 133788 4626 133840 4632
rect 133800 2990 133828 4626
rect 133788 2984 133840 2990
rect 133788 2926 133840 2932
rect 132960 2168 133012 2174
rect 132960 2110 133012 2116
rect 132972 480 133000 2110
rect 133788 1488 133840 1494
rect 133788 1430 133840 1436
rect 133800 1018 133828 1430
rect 133788 1012 133840 1018
rect 133788 954 133840 960
rect 134168 480 134196 6870
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 135076 2168 135128 2174
rect 135076 2110 135128 2116
rect 135088 1057 135116 2110
rect 135074 1048 135130 1057
rect 135074 983 135130 992
rect 135272 480 135300 3334
rect 136272 1420 136324 1426
rect 136272 1362 136324 1368
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136284 474 136312 1362
rect 136468 480 136496 6886
rect 137940 4622 137968 8230
rect 139320 6914 139348 8774
rect 139320 6886 139532 6914
rect 139400 4752 139452 4758
rect 139400 4694 139452 4700
rect 137928 4616 137980 4622
rect 137928 4558 137980 4564
rect 137652 4072 137704 4078
rect 137652 4014 137704 4020
rect 137284 1692 137336 1698
rect 137284 1634 137336 1640
rect 136548 1556 136600 1562
rect 136548 1498 136600 1504
rect 136560 1329 136588 1498
rect 137296 1358 137324 1634
rect 137284 1352 137336 1358
rect 136546 1320 136602 1329
rect 137284 1294 137336 1300
rect 136546 1255 136602 1264
rect 137664 480 137692 4014
rect 139412 2990 139440 4694
rect 138848 2984 138900 2990
rect 138848 2926 138900 2932
rect 139400 2984 139452 2990
rect 139400 2926 139452 2932
rect 138860 480 138888 2926
rect 139504 1222 139532 6886
rect 140148 5914 140176 12514
rect 140780 10056 140832 10062
rect 140780 9998 140832 10004
rect 140792 8809 140820 9998
rect 143092 9654 143120 15642
rect 143080 9648 143132 9654
rect 143080 9590 143132 9596
rect 143908 9648 143960 9654
rect 143908 9590 143960 9596
rect 140778 8800 140834 8809
rect 140778 8735 140834 8744
rect 143540 7540 143592 7546
rect 143540 7482 143592 7488
rect 140780 7404 140832 7410
rect 140780 7346 140832 7352
rect 140686 6080 140742 6089
rect 140686 6015 140742 6024
rect 140700 5982 140728 6015
rect 140688 5976 140740 5982
rect 140688 5918 140740 5924
rect 140136 5908 140188 5914
rect 140136 5850 140188 5856
rect 140792 2038 140820 7346
rect 143552 5681 143580 7482
rect 143538 5672 143594 5681
rect 143538 5607 143594 5616
rect 142436 2984 142488 2990
rect 142436 2926 142488 2932
rect 141240 2916 141292 2922
rect 141240 2858 141292 2864
rect 140780 2032 140832 2038
rect 140780 1974 140832 1980
rect 140044 1488 140096 1494
rect 140044 1430 140096 1436
rect 139492 1216 139544 1222
rect 139492 1158 139544 1164
rect 140056 480 140084 1430
rect 141252 480 141280 2858
rect 142448 480 142476 2926
rect 143920 2650 143948 9590
rect 144644 6044 144696 6050
rect 144644 5986 144696 5992
rect 145012 6044 145064 6050
rect 145012 5986 145064 5992
rect 143908 2644 143960 2650
rect 143908 2586 143960 2592
rect 142804 1624 142856 1630
rect 142804 1566 142856 1572
rect 142816 1018 142844 1566
rect 144656 1442 144684 5986
rect 144736 5500 144788 5506
rect 144736 5442 144788 5448
rect 144748 2854 144776 5442
rect 144828 4276 144880 4282
rect 144828 4218 144880 4224
rect 144736 2848 144788 2854
rect 144736 2790 144788 2796
rect 144840 2174 144868 4218
rect 145024 2417 145052 5986
rect 146668 5908 146720 5914
rect 146668 5850 146720 5856
rect 146576 4752 146628 4758
rect 146576 4694 146628 4700
rect 145932 4140 145984 4146
rect 145932 4082 145984 4088
rect 145010 2408 145066 2417
rect 145010 2343 145066 2352
rect 144828 2168 144880 2174
rect 144828 2110 144880 2116
rect 144920 2168 144972 2174
rect 144920 2110 144972 2116
rect 142896 1420 142948 1426
rect 144656 1414 144776 1442
rect 142896 1362 142948 1368
rect 142804 1012 142856 1018
rect 142804 954 142856 960
rect 142908 950 142936 1362
rect 142896 944 142948 950
rect 142896 886 142948 892
rect 144748 480 144776 1414
rect 144932 814 144960 2110
rect 144920 808 144972 814
rect 144920 750 144972 756
rect 145944 480 145972 4082
rect 146588 2553 146616 4694
rect 146680 3330 146708 5850
rect 146864 3482 146892 16546
rect 146956 8294 146984 18498
rect 147692 17921 147720 18974
rect 147772 18148 147824 18154
rect 147772 18090 147824 18096
rect 147678 17912 147734 17921
rect 147678 17847 147734 17856
rect 147784 17762 147812 18090
rect 147692 17734 147812 17762
rect 147692 16590 147720 17734
rect 147680 16584 147732 16590
rect 147680 16526 147732 16532
rect 148336 12442 148364 19450
rect 149072 19174 149100 19654
rect 150440 19644 150492 19650
rect 150440 19586 150492 19592
rect 150452 19242 150480 19586
rect 150440 19236 150492 19242
rect 150440 19178 150492 19184
rect 149060 19168 149112 19174
rect 149060 19110 149112 19116
rect 149244 19032 149296 19038
rect 149244 18974 149296 18980
rect 149152 18556 149204 18562
rect 149152 18498 149204 18504
rect 149060 18352 149112 18358
rect 149060 18294 149112 18300
rect 149072 17882 149100 18294
rect 149060 17876 149112 17882
rect 149060 17818 149112 17824
rect 149164 17066 149192 18498
rect 149152 17060 149204 17066
rect 149152 17002 149204 17008
rect 149256 16574 149284 18974
rect 150532 18488 150584 18494
rect 150532 18430 150584 18436
rect 148980 16546 149284 16574
rect 148980 14142 149008 16546
rect 150440 15836 150492 15842
rect 150440 15778 150492 15784
rect 150452 15094 150480 15778
rect 150440 15088 150492 15094
rect 150440 15030 150492 15036
rect 148968 14136 149020 14142
rect 148968 14078 149020 14084
rect 149060 13864 149112 13870
rect 149060 13806 149112 13812
rect 148324 12436 148376 12442
rect 148324 12378 148376 12384
rect 149072 11393 149100 13806
rect 150544 13569 150572 18430
rect 150636 18154 150664 19790
rect 150624 18148 150676 18154
rect 150624 18090 150676 18096
rect 150530 13560 150586 13569
rect 150530 13495 150586 13504
rect 149058 11384 149114 11393
rect 149058 11319 149114 11328
rect 147036 10260 147088 10266
rect 147036 10202 147088 10208
rect 146944 8288 146996 8294
rect 146944 8230 146996 8236
rect 147048 6089 147076 10202
rect 149612 8288 149664 8294
rect 149612 8230 149664 8236
rect 149244 8220 149296 8226
rect 149244 8162 149296 8168
rect 147034 6080 147090 6089
rect 147034 6015 147090 6024
rect 149152 5500 149204 5506
rect 149152 5442 149204 5448
rect 149164 4758 149192 5442
rect 149152 4752 149204 4758
rect 146942 4720 146998 4729
rect 149152 4694 149204 4700
rect 146942 4655 146998 4664
rect 146956 4078 146984 4655
rect 146944 4072 146996 4078
rect 146944 4014 146996 4020
rect 146864 3454 147168 3482
rect 146668 3324 146720 3330
rect 146668 3266 146720 3272
rect 146574 2544 146630 2553
rect 146574 2479 146630 2488
rect 146300 1556 146352 1562
rect 146300 1498 146352 1504
rect 146312 1290 146340 1498
rect 146300 1284 146352 1290
rect 146300 1226 146352 1232
rect 147140 480 147168 3454
rect 149060 1488 149112 1494
rect 149060 1430 149112 1436
rect 148324 1352 148376 1358
rect 148324 1294 148376 1300
rect 148336 480 148364 1294
rect 136272 468 136324 474
rect 136272 410 136324 416
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 82 143622 480
rect 143368 66 143622 82
rect 143356 60 143622 66
rect 143408 54 143622 60
rect 143356 2 143408 8
rect 143510 -960 143622 54
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149072 270 149100 1430
rect 149256 1290 149284 8162
rect 149520 3392 149572 3398
rect 149520 3334 149572 3340
rect 149244 1284 149296 1290
rect 149244 1226 149296 1232
rect 149532 480 149560 3334
rect 149624 2786 149652 8230
rect 150532 6996 150584 7002
rect 150532 6938 150584 6944
rect 150440 6928 150492 6934
rect 150440 6870 150492 6876
rect 150452 6118 150480 6870
rect 150440 6112 150492 6118
rect 150440 6054 150492 6060
rect 150440 5568 150492 5574
rect 150440 5510 150492 5516
rect 150452 4049 150480 5510
rect 150544 4282 150572 6938
rect 150728 6914 150756 160890
rect 150808 159588 150860 159594
rect 150808 159530 150860 159536
rect 150636 6886 150756 6914
rect 150532 4276 150584 4282
rect 150532 4218 150584 4224
rect 150438 4040 150494 4049
rect 150438 3975 150494 3984
rect 150440 3052 150492 3058
rect 150440 2994 150492 3000
rect 149612 2780 149664 2786
rect 149612 2722 149664 2728
rect 150452 1834 150480 2994
rect 150440 1828 150492 1834
rect 150440 1770 150492 1776
rect 150636 480 150664 6886
rect 150820 1358 150848 159530
rect 151176 155372 151228 155378
rect 151176 155314 151228 155320
rect 151082 155272 151138 155281
rect 151082 155207 151138 155216
rect 150992 152516 151044 152522
rect 150992 152458 151044 152464
rect 150898 151872 150954 151881
rect 150898 151807 150954 151816
rect 150912 151638 150940 151807
rect 150900 151632 150952 151638
rect 150900 151574 150952 151580
rect 151004 151094 151032 152458
rect 150992 151088 151044 151094
rect 150992 151030 151044 151036
rect 151096 100706 151124 155207
rect 151188 139398 151216 155314
rect 151452 154692 151504 154698
rect 151452 154634 151504 154640
rect 151360 154012 151412 154018
rect 151360 153954 151412 153960
rect 151266 153368 151322 153377
rect 151266 153303 151322 153312
rect 151280 151162 151308 153303
rect 151372 151434 151400 153954
rect 151360 151428 151412 151434
rect 151360 151370 151412 151376
rect 151464 151230 151492 154634
rect 151452 151224 151504 151230
rect 151452 151166 151504 151172
rect 151268 151156 151320 151162
rect 151268 151098 151320 151104
rect 151176 139392 151228 139398
rect 151176 139334 151228 139340
rect 151084 100700 151136 100706
rect 151084 100642 151136 100648
rect 150900 22908 150952 22914
rect 150900 22850 150952 22856
rect 150912 19922 150940 22850
rect 151360 22704 151412 22710
rect 151360 22646 151412 22652
rect 150992 22160 151044 22166
rect 150992 22102 151044 22108
rect 150900 19916 150952 19922
rect 150900 19858 150952 19864
rect 151004 19689 151032 22102
rect 151268 20664 151320 20670
rect 151268 20606 151320 20612
rect 151084 19984 151136 19990
rect 151084 19926 151136 19932
rect 150990 19680 151046 19689
rect 150990 19615 151046 19624
rect 151096 19106 151124 19926
rect 151176 19780 151228 19786
rect 151176 19722 151228 19728
rect 151084 19100 151136 19106
rect 151084 19042 151136 19048
rect 151188 18170 151216 19722
rect 151280 19038 151308 20606
rect 151268 19032 151320 19038
rect 151268 18974 151320 18980
rect 151268 18896 151320 18902
rect 151268 18838 151320 18844
rect 150900 18148 150952 18154
rect 150900 18090 150952 18096
rect 151096 18142 151216 18170
rect 150912 12209 150940 18090
rect 150898 12200 150954 12209
rect 150898 12135 150954 12144
rect 151096 5642 151124 18142
rect 151176 18012 151228 18018
rect 151176 17954 151228 17960
rect 151188 9489 151216 17954
rect 151174 9480 151230 9489
rect 151174 9415 151230 9424
rect 151280 8226 151308 18838
rect 151372 11422 151400 22646
rect 151452 21072 151504 21078
rect 151452 21014 151504 21020
rect 151464 18018 151492 21014
rect 151544 20324 151596 20330
rect 151544 20266 151596 20272
rect 151452 18012 151504 18018
rect 151452 17954 151504 17960
rect 151556 17202 151584 20266
rect 151544 17196 151596 17202
rect 151544 17138 151596 17144
rect 151360 11416 151412 11422
rect 151360 11358 151412 11364
rect 151832 11014 151860 162250
rect 153844 162240 153896 162246
rect 153844 162182 153896 162188
rect 152648 160880 152700 160886
rect 152648 160822 152700 160828
rect 152464 159520 152516 159526
rect 152464 159462 152516 159468
rect 151912 158092 151964 158098
rect 151912 158034 151964 158040
rect 151924 18562 151952 158034
rect 152094 153232 152150 153241
rect 152094 153167 152150 153176
rect 152004 152720 152056 152726
rect 152004 152662 152056 152668
rect 152016 151366 152044 152662
rect 152004 151360 152056 151366
rect 152004 151302 152056 151308
rect 152108 151298 152136 153167
rect 152096 151292 152148 151298
rect 152096 151234 152148 151240
rect 152476 32434 152504 159462
rect 152554 153776 152610 153785
rect 152554 153711 152610 153720
rect 152568 46918 152596 153711
rect 152660 75886 152688 160822
rect 152740 156596 152792 156602
rect 152740 156538 152792 156544
rect 152752 149734 152780 156538
rect 153108 155236 153160 155242
rect 153108 155178 153160 155184
rect 152924 154760 152976 154766
rect 152924 154702 152976 154708
rect 152832 154692 152884 154698
rect 152832 154634 152884 154640
rect 152844 151502 152872 154634
rect 152936 151570 152964 154702
rect 153120 154154 153148 155178
rect 153108 154148 153160 154154
rect 153108 154090 153160 154096
rect 152924 151564 152976 151570
rect 152924 151506 152976 151512
rect 152832 151496 152884 151502
rect 152832 151438 152884 151444
rect 152740 149728 152792 149734
rect 152740 149670 152792 149676
rect 152648 75880 152700 75886
rect 152648 75822 152700 75828
rect 152556 46912 152608 46918
rect 152556 46854 152608 46860
rect 152464 32428 152516 32434
rect 152464 32370 152516 32376
rect 153856 31142 153884 162182
rect 156604 159656 156656 159662
rect 156604 159598 156656 159604
rect 155868 158228 155920 158234
rect 155868 158170 155920 158176
rect 154028 158024 154080 158030
rect 154028 157966 154080 157972
rect 153934 153912 153990 153921
rect 153934 153847 153990 153856
rect 153948 86970 153976 153847
rect 154040 149802 154068 157966
rect 154120 155576 154172 155582
rect 154120 155518 154172 155524
rect 154132 149870 154160 155518
rect 155880 155242 155908 158170
rect 156512 155440 156564 155446
rect 156512 155382 156564 155388
rect 155868 155236 155920 155242
rect 155868 155178 155920 155184
rect 156524 153950 156552 155382
rect 156616 154018 156644 159598
rect 161480 159452 161532 159458
rect 161480 159394 161532 159400
rect 160100 156528 160152 156534
rect 160100 156470 160152 156476
rect 156696 155304 156748 155310
rect 156696 155246 156748 155252
rect 156604 154012 156656 154018
rect 156604 153954 156656 153960
rect 156512 153944 156564 153950
rect 156512 153886 156564 153892
rect 156604 153672 156656 153678
rect 156604 153614 156656 153620
rect 154120 149864 154172 149870
rect 154120 149806 154172 149812
rect 154028 149796 154080 149802
rect 154028 149738 154080 149744
rect 153936 86964 153988 86970
rect 153936 86906 153988 86912
rect 156616 74390 156644 153614
rect 156708 152522 156736 155246
rect 160112 154086 160140 156470
rect 160100 154080 160152 154086
rect 160100 154022 160152 154028
rect 157982 153504 158038 153513
rect 157982 153439 158038 153448
rect 156696 152516 156748 152522
rect 156696 152458 156748 152464
rect 156694 152416 156750 152425
rect 156694 152351 156750 152360
rect 156708 126954 156736 152351
rect 156696 126948 156748 126954
rect 156696 126890 156748 126896
rect 156696 75880 156748 75886
rect 156696 75822 156748 75828
rect 156604 74384 156656 74390
rect 156604 74326 156656 74332
rect 153844 31136 153896 31142
rect 153844 31078 153896 31084
rect 156708 31074 156736 75822
rect 157996 33114 158024 153439
rect 160742 152280 160798 152289
rect 160742 152215 160798 152224
rect 160100 74384 160152 74390
rect 160100 74326 160152 74332
rect 157984 33108 158036 33114
rect 157984 33050 158036 33056
rect 156696 31068 156748 31074
rect 156696 31010 156748 31016
rect 153292 26716 153344 26722
rect 153292 26658 153344 26664
rect 152096 26580 152148 26586
rect 152096 26522 152148 26528
rect 152108 22914 152136 26522
rect 152924 25084 152976 25090
rect 152924 25026 152976 25032
rect 152832 23792 152884 23798
rect 152832 23734 152884 23740
rect 152648 23452 152700 23458
rect 152648 23394 152700 23400
rect 152096 22908 152148 22914
rect 152096 22850 152148 22856
rect 152556 21004 152608 21010
rect 152556 20946 152608 20952
rect 152004 20936 152056 20942
rect 152004 20878 152056 20884
rect 151912 18556 151964 18562
rect 151912 18498 151964 18504
rect 152016 18034 152044 20878
rect 152372 20664 152424 20670
rect 152372 20606 152424 20612
rect 152188 19576 152240 19582
rect 152188 19518 152240 19524
rect 152200 18154 152228 19518
rect 152188 18148 152240 18154
rect 152188 18090 152240 18096
rect 151924 18006 152044 18034
rect 151924 17950 151952 18006
rect 151912 17944 151964 17950
rect 151912 17886 151964 17892
rect 152004 17944 152056 17950
rect 152004 17886 152056 17892
rect 152016 15434 152044 17886
rect 152004 15428 152056 15434
rect 152004 15370 152056 15376
rect 151360 11008 151412 11014
rect 151360 10950 151412 10956
rect 151820 11008 151872 11014
rect 151820 10950 151872 10956
rect 151268 8220 151320 8226
rect 151268 8162 151320 8168
rect 151084 5636 151136 5642
rect 151084 5578 151136 5584
rect 151372 3398 151400 10950
rect 152384 7546 152412 20606
rect 152464 19916 152516 19922
rect 152464 19858 152516 19864
rect 152476 19718 152504 19858
rect 152568 19854 152596 20946
rect 152556 19848 152608 19854
rect 152556 19790 152608 19796
rect 152464 19712 152516 19718
rect 152464 19654 152516 19660
rect 152556 19712 152608 19718
rect 152556 19654 152608 19660
rect 152568 9625 152596 19654
rect 152660 16561 152688 23394
rect 152740 20052 152792 20058
rect 152740 19994 152792 20000
rect 152646 16552 152702 16561
rect 152646 16487 152702 16496
rect 152752 13870 152780 19994
rect 152844 18970 152872 23734
rect 152936 20330 152964 25026
rect 153108 24880 153160 24886
rect 153108 24822 153160 24828
rect 153016 22432 153068 22438
rect 153016 22374 153068 22380
rect 152924 20324 152976 20330
rect 152924 20266 152976 20272
rect 153028 19786 153056 22374
rect 153120 22166 153148 24822
rect 153108 22160 153160 22166
rect 153108 22102 153160 22108
rect 153304 20738 153332 26658
rect 157248 26648 157300 26654
rect 157248 26590 157300 26596
rect 156972 26376 157024 26382
rect 156972 26318 157024 26324
rect 154948 26308 155000 26314
rect 154948 26250 155000 26256
rect 153384 25288 153436 25294
rect 153384 25230 153436 25236
rect 153292 20732 153344 20738
rect 153292 20674 153344 20680
rect 153292 20596 153344 20602
rect 153292 20538 153344 20544
rect 153108 20120 153160 20126
rect 153108 20062 153160 20068
rect 153016 19780 153068 19786
rect 153016 19722 153068 19728
rect 152832 18964 152884 18970
rect 152832 18906 152884 18912
rect 153016 18284 153068 18290
rect 153016 18226 153068 18232
rect 153028 17921 153056 18226
rect 153014 17912 153070 17921
rect 153014 17847 153070 17856
rect 153120 17649 153148 20062
rect 153304 19281 153332 20538
rect 153396 19922 153424 25230
rect 154028 22568 154080 22574
rect 154028 22510 154080 22516
rect 153936 22228 153988 22234
rect 153936 22170 153988 22176
rect 153844 21276 153896 21282
rect 153844 21218 153896 21224
rect 153384 19916 153436 19922
rect 153384 19858 153436 19864
rect 153752 19848 153804 19854
rect 153752 19790 153804 19796
rect 153660 19304 153712 19310
rect 153290 19272 153346 19281
rect 153660 19246 153712 19252
rect 153290 19207 153346 19216
rect 153106 17640 153162 17649
rect 153106 17575 153162 17584
rect 153672 16658 153700 19246
rect 153660 16652 153712 16658
rect 153660 16594 153712 16600
rect 153108 15768 153160 15774
rect 153108 15710 153160 15716
rect 153120 15298 153148 15710
rect 153764 15609 153792 19790
rect 153750 15600 153806 15609
rect 153750 15535 153806 15544
rect 153108 15292 153160 15298
rect 153108 15234 153160 15240
rect 152740 13864 152792 13870
rect 152740 13806 152792 13812
rect 152554 9616 152610 9625
rect 152554 9551 152610 9560
rect 152372 7540 152424 7546
rect 152372 7482 152424 7488
rect 153752 4412 153804 4418
rect 153752 4354 153804 4360
rect 152924 3936 152976 3942
rect 152924 3878 152976 3884
rect 151360 3392 151412 3398
rect 151360 3334 151412 3340
rect 151820 1964 151872 1970
rect 151820 1906 151872 1912
rect 150808 1352 150860 1358
rect 150808 1294 150860 1300
rect 151832 480 151860 1906
rect 152936 1034 152964 3878
rect 153016 2848 153068 2854
rect 153016 2790 153068 2796
rect 153028 1222 153056 2790
rect 153764 2650 153792 4354
rect 153856 3058 153884 21218
rect 153948 16833 153976 22170
rect 154040 18873 154068 22510
rect 154212 22500 154264 22506
rect 154212 22442 154264 22448
rect 154120 20800 154172 20806
rect 154120 20742 154172 20748
rect 154026 18864 154082 18873
rect 154026 18799 154082 18808
rect 154132 18714 154160 20742
rect 154224 19650 154252 22442
rect 154304 22296 154356 22302
rect 154304 22238 154356 22244
rect 154212 19644 154264 19650
rect 154212 19586 154264 19592
rect 154316 19530 154344 22238
rect 154396 21208 154448 21214
rect 154396 21150 154448 21156
rect 154040 18686 154160 18714
rect 154224 19502 154344 19530
rect 153934 16824 153990 16833
rect 153934 16759 153990 16768
rect 153936 16652 153988 16658
rect 153936 16594 153988 16600
rect 153948 7002 153976 16594
rect 154040 10266 154068 18686
rect 154224 18578 154252 19502
rect 154304 19236 154356 19242
rect 154304 19178 154356 19184
rect 154132 18550 154252 18578
rect 154132 11529 154160 18550
rect 154212 18148 154264 18154
rect 154212 18090 154264 18096
rect 154118 11520 154174 11529
rect 154118 11455 154174 11464
rect 154028 10260 154080 10266
rect 154028 10202 154080 10208
rect 154224 9058 154252 18090
rect 154316 13433 154344 19178
rect 154408 15201 154436 21150
rect 154488 20868 154540 20874
rect 154488 20810 154540 20816
rect 154500 18494 154528 20810
rect 154960 20602 154988 26250
rect 156052 25220 156104 25226
rect 156052 25162 156104 25168
rect 155776 23860 155828 23866
rect 155776 23802 155828 23808
rect 155132 23520 155184 23526
rect 155132 23462 155184 23468
rect 155144 20942 155172 23462
rect 155684 21344 155736 21350
rect 155684 21286 155736 21292
rect 155132 20936 155184 20942
rect 155132 20878 155184 20884
rect 155224 20936 155276 20942
rect 155224 20878 155276 20884
rect 154948 20596 155000 20602
rect 154948 20538 155000 20544
rect 154580 19508 154632 19514
rect 154580 19450 154632 19456
rect 154592 19242 154620 19450
rect 154580 19236 154632 19242
rect 154580 19178 154632 19184
rect 154488 18488 154540 18494
rect 154488 18430 154540 18436
rect 154394 15192 154450 15201
rect 154394 15127 154450 15136
rect 154302 13424 154358 13433
rect 154302 13359 154358 13368
rect 154304 9580 154356 9586
rect 154304 9522 154356 9528
rect 154132 9030 154252 9058
rect 154132 8809 154160 9030
rect 154212 8900 154264 8906
rect 154212 8842 154264 8848
rect 154118 8800 154174 8809
rect 154118 8735 154174 8744
rect 153936 6996 153988 7002
rect 153936 6938 153988 6944
rect 153844 3052 153896 3058
rect 153844 2994 153896 3000
rect 153752 2644 153804 2650
rect 153752 2586 153804 2592
rect 153108 2100 153160 2106
rect 153108 2042 153160 2048
rect 153016 1216 153068 1222
rect 153016 1158 153068 1164
rect 152936 1006 153056 1034
rect 153028 480 153056 1006
rect 153120 882 153148 2042
rect 153108 876 153160 882
rect 153108 818 153160 824
rect 154224 480 154252 8842
rect 154316 5574 154344 9522
rect 154304 5568 154356 5574
rect 154304 5510 154356 5516
rect 155236 5506 155264 20878
rect 155500 20188 155552 20194
rect 155500 20130 155552 20136
rect 155316 19780 155368 19786
rect 155316 19722 155368 19728
rect 155328 8158 155356 19722
rect 155408 15224 155460 15230
rect 155408 15166 155460 15172
rect 155316 8152 155368 8158
rect 155316 8094 155368 8100
rect 155420 6050 155448 15166
rect 155512 13705 155540 20130
rect 155696 16425 155724 21286
rect 155788 18902 155816 23802
rect 155960 21412 156012 21418
rect 155960 21354 156012 21360
rect 155868 21140 155920 21146
rect 155868 21082 155920 21088
rect 155880 19990 155908 21082
rect 155868 19984 155920 19990
rect 155868 19926 155920 19932
rect 155972 19802 156000 21354
rect 155880 19774 156000 19802
rect 155776 18896 155828 18902
rect 155776 18838 155828 18844
rect 155880 18154 155908 19774
rect 155960 19644 156012 19650
rect 155960 19586 156012 19592
rect 155868 18148 155920 18154
rect 155868 18090 155920 18096
rect 155972 16574 156000 19586
rect 156064 19310 156092 25162
rect 156604 25152 156656 25158
rect 156604 25094 156656 25100
rect 156512 22364 156564 22370
rect 156512 22306 156564 22312
rect 156524 19854 156552 22306
rect 156616 20126 156644 25094
rect 156696 23656 156748 23662
rect 156696 23598 156748 23604
rect 156604 20120 156656 20126
rect 156604 20062 156656 20068
rect 156512 19848 156564 19854
rect 156512 19790 156564 19796
rect 156604 19848 156656 19854
rect 156604 19790 156656 19796
rect 156052 19304 156104 19310
rect 156052 19246 156104 19252
rect 155880 16546 156000 16574
rect 155682 16416 155738 16425
rect 155682 16351 155738 16360
rect 155498 13696 155554 13705
rect 155498 13631 155554 13640
rect 155880 12442 155908 16546
rect 155960 13796 156012 13802
rect 155960 13738 156012 13744
rect 155868 12436 155920 12442
rect 155868 12378 155920 12384
rect 155972 12073 156000 13738
rect 155958 12064 156014 12073
rect 155958 11999 156014 12008
rect 156512 9784 156564 9790
rect 156512 9726 156564 9732
rect 156524 7070 156552 9726
rect 156512 7064 156564 7070
rect 156512 7006 156564 7012
rect 155408 6044 155460 6050
rect 155408 5986 155460 5992
rect 155224 5500 155276 5506
rect 155224 5442 155276 5448
rect 156616 4418 156644 19790
rect 156708 10985 156736 23598
rect 156984 20194 157012 26318
rect 157064 23588 157116 23594
rect 157064 23530 157116 23536
rect 157076 21350 157104 23530
rect 157064 21344 157116 21350
rect 157064 21286 157116 21292
rect 157260 20942 157288 26590
rect 159364 26512 159416 26518
rect 159364 26454 159416 26460
rect 157340 26444 157392 26450
rect 157340 26386 157392 26392
rect 157248 20936 157300 20942
rect 157248 20878 157300 20884
rect 157352 20754 157380 26386
rect 157892 25016 157944 25022
rect 157892 24958 157944 24964
rect 157432 22636 157484 22642
rect 157432 22578 157484 22584
rect 157260 20726 157380 20754
rect 156972 20188 157024 20194
rect 156972 20130 157024 20136
rect 156788 19916 156840 19922
rect 156788 19858 156840 19864
rect 156800 12986 156828 19858
rect 157260 19718 157288 20726
rect 157248 19712 157300 19718
rect 157248 19654 157300 19660
rect 157444 18426 157472 22578
rect 157904 21418 157932 24958
rect 158076 23928 158128 23934
rect 158076 23870 158128 23876
rect 157892 21412 157944 21418
rect 157892 21354 157944 21360
rect 157984 20732 158036 20738
rect 157984 20674 158036 20680
rect 157800 20052 157852 20058
rect 157800 19994 157852 20000
rect 157708 19780 157760 19786
rect 157708 19722 157760 19728
rect 157720 19514 157748 19722
rect 157812 19514 157840 19994
rect 157708 19508 157760 19514
rect 157708 19450 157760 19456
rect 157800 19508 157852 19514
rect 157800 19450 157852 19456
rect 157432 18420 157484 18426
rect 157432 18362 157484 18368
rect 157340 14068 157392 14074
rect 157340 14010 157392 14016
rect 156788 12980 156840 12986
rect 156788 12922 156840 12928
rect 157352 12753 157380 14010
rect 157338 12744 157394 12753
rect 157338 12679 157394 12688
rect 156694 10976 156750 10985
rect 156694 10911 156750 10920
rect 156972 9648 157024 9654
rect 156972 9590 157024 9596
rect 156604 4412 156656 4418
rect 156604 4354 156656 4360
rect 156604 4004 156656 4010
rect 156604 3946 156656 3952
rect 155408 3392 155460 3398
rect 155408 3334 155460 3340
rect 154488 2916 154540 2922
rect 154488 2858 154540 2864
rect 154500 2038 154528 2858
rect 154488 2032 154540 2038
rect 154488 1974 154540 1980
rect 155420 480 155448 3334
rect 156616 480 156644 3946
rect 156984 3194 157012 9590
rect 157996 4078 158024 20674
rect 158088 9586 158116 23870
rect 158168 22160 158220 22166
rect 158168 22102 158220 22108
rect 158180 15842 158208 22102
rect 158260 21344 158312 21350
rect 158260 21286 158312 21292
rect 158272 16590 158300 21286
rect 158444 18148 158496 18154
rect 158444 18090 158496 18096
rect 158260 16584 158312 16590
rect 158260 16526 158312 16532
rect 158168 15836 158220 15842
rect 158168 15778 158220 15784
rect 158456 15162 158484 18090
rect 158444 15156 158496 15162
rect 158444 15098 158496 15104
rect 159376 9654 159404 26454
rect 159456 24948 159508 24954
rect 159456 24890 159508 24896
rect 159468 13802 159496 24890
rect 159548 23996 159600 24002
rect 159548 23938 159600 23944
rect 159560 14074 159588 23938
rect 159548 14068 159600 14074
rect 159548 14010 159600 14016
rect 159456 13796 159508 13802
rect 159456 13738 159508 13744
rect 159364 9648 159416 9654
rect 159364 9590 159416 9596
rect 158076 9580 158128 9586
rect 158076 9522 158128 9528
rect 157984 4072 158036 4078
rect 157984 4014 158036 4020
rect 160112 3398 160140 74326
rect 160756 73166 160784 152215
rect 160744 73160 160796 73166
rect 160744 73102 160796 73108
rect 160192 25356 160244 25362
rect 160192 25298 160244 25304
rect 160204 21350 160232 25298
rect 160192 21344 160244 21350
rect 160192 21286 160244 21292
rect 160192 18012 160244 18018
rect 160192 17954 160244 17960
rect 160204 17202 160232 17954
rect 160192 17196 160244 17202
rect 160192 17138 160244 17144
rect 161492 16574 161520 159394
rect 169772 159361 169800 702406
rect 201512 171834 201540 702986
rect 218992 699718 219020 703520
rect 217324 699712 217376 699718
rect 217324 699654 217376 699660
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 217336 173194 217364 699654
rect 234632 494766 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 693462 267688 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 267648 693456 267700 693462
rect 267648 693398 267700 693404
rect 234620 494760 234672 494766
rect 234620 494702 234672 494708
rect 217324 173188 217376 173194
rect 217324 173130 217376 173136
rect 201500 171828 201552 171834
rect 201500 171770 201552 171776
rect 188344 162172 188396 162178
rect 188344 162114 188396 162120
rect 174544 160812 174596 160818
rect 174544 160754 174596 160760
rect 169758 159352 169814 159361
rect 169758 159287 169814 159296
rect 163502 157448 163558 157457
rect 163502 157383 163558 157392
rect 163516 155310 163544 157383
rect 164240 155780 164292 155786
rect 164240 155722 164292 155728
rect 163504 155304 163556 155310
rect 163504 155246 163556 155252
rect 162122 153640 162178 153649
rect 162122 153575 162178 153584
rect 162136 113150 162164 153575
rect 162124 113144 162176 113150
rect 162124 113086 162176 113092
rect 164252 16574 164280 155722
rect 171140 154828 171192 154834
rect 171140 154770 171192 154776
rect 164792 154148 164844 154154
rect 164792 154090 164844 154096
rect 164804 152726 164832 154090
rect 164792 152720 164844 152726
rect 164792 152662 164844 152668
rect 166264 152652 166316 152658
rect 166264 152594 166316 152600
rect 165896 32428 165948 32434
rect 165896 32370 165948 32376
rect 165908 30326 165936 32370
rect 166276 31414 166304 152594
rect 166264 31408 166316 31414
rect 166264 31350 166316 31356
rect 168472 31408 168524 31414
rect 168472 31350 168524 31356
rect 165896 30320 165948 30326
rect 165896 30262 165948 30268
rect 161492 16546 162072 16574
rect 164252 16546 164464 16574
rect 160192 12300 160244 12306
rect 160192 12242 160244 12248
rect 160204 8906 160232 12242
rect 160192 8900 160244 8906
rect 160192 8842 160244 8848
rect 160560 6928 160612 6934
rect 160560 6870 160612 6876
rect 160190 3768 160246 3777
rect 160190 3703 160246 3712
rect 160100 3392 160152 3398
rect 160100 3334 160152 3340
rect 156972 3188 157024 3194
rect 156972 3130 157024 3136
rect 157340 3052 157392 3058
rect 157340 2994 157392 3000
rect 157352 2514 157380 2994
rect 157800 2916 157852 2922
rect 157800 2858 157852 2864
rect 157340 2508 157392 2514
rect 157340 2450 157392 2456
rect 157812 480 157840 2858
rect 158904 2848 158956 2854
rect 158904 2790 158956 2796
rect 158812 2440 158864 2446
rect 158812 2382 158864 2388
rect 158720 1420 158772 1426
rect 158720 1362 158772 1368
rect 149060 264 149112 270
rect 149060 206 149112 212
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158732 202 158760 1362
rect 158824 1018 158852 2382
rect 158812 1012 158864 1018
rect 158812 954 158864 960
rect 158916 480 158944 2790
rect 160204 1442 160232 3703
rect 160572 3330 160600 6870
rect 161296 3392 161348 3398
rect 161296 3334 161348 3340
rect 160560 3324 160612 3330
rect 160560 3266 160612 3272
rect 160112 1414 160232 1442
rect 160112 480 160140 1414
rect 161308 480 161336 3334
rect 158720 196 158772 202
rect 158720 138 158772 144
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 162860 8628 162912 8634
rect 162860 8570 162912 8576
rect 162872 3194 162900 8570
rect 163688 3324 163740 3330
rect 163688 3266 163740 3272
rect 162860 3188 162912 3194
rect 162860 3130 162912 3136
rect 163700 480 163728 3266
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 167184 15360 167236 15366
rect 167184 15302 167236 15308
rect 166080 9988 166132 9994
rect 166080 9930 166132 9936
rect 166092 480 166120 9930
rect 167196 480 167224 15302
rect 168380 13048 168432 13054
rect 168380 12990 168432 12996
rect 168392 12442 168420 12990
rect 168380 12436 168432 12442
rect 168380 12378 168432 12384
rect 168484 6914 168512 31350
rect 171152 16574 171180 154770
rect 172520 30320 172572 30326
rect 172520 30262 172572 30268
rect 172532 16574 172560 30262
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 168564 14204 168616 14210
rect 168564 14146 168616 14152
rect 168576 12986 168604 14146
rect 168564 12980 168616 12986
rect 168564 12922 168616 12928
rect 170312 12368 170364 12374
rect 170312 12310 170364 12316
rect 168392 6886 168512 6914
rect 168392 480 168420 6886
rect 169576 3188 169628 3194
rect 169576 3130 169628 3136
rect 169588 480 169616 3130
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 12310
rect 171980 480 172008 16546
rect 172520 8560 172572 8566
rect 172520 8502 172572 8508
rect 172532 3942 172560 8502
rect 172520 3936 172572 3942
rect 172520 3878 172572 3884
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 174268 5840 174320 5846
rect 174268 5782 174320 5788
rect 173532 2508 173584 2514
rect 173532 2450 173584 2456
rect 173544 1086 173572 2450
rect 173532 1080 173584 1086
rect 173532 1022 173584 1028
rect 174280 480 174308 5782
rect 174556 3398 174584 160754
rect 180064 159384 180116 159390
rect 180064 159326 180116 159332
rect 175280 152720 175332 152726
rect 175280 152662 175332 152668
rect 175292 16574 175320 152662
rect 178040 152584 178092 152590
rect 178040 152526 178092 152532
rect 176752 22704 176804 22710
rect 176752 22646 176804 22652
rect 176764 16574 176792 22646
rect 178052 16574 178080 152526
rect 179420 31136 179472 31142
rect 179420 31078 179472 31084
rect 178132 19916 178184 19922
rect 178132 19858 178184 19864
rect 178144 18902 178172 19858
rect 178132 18896 178184 18902
rect 178132 18838 178184 18844
rect 179432 16574 179460 31078
rect 180076 29646 180104 159326
rect 184940 154896 184992 154902
rect 184940 154838 184992 154844
rect 182180 151632 182232 151638
rect 182180 151574 182232 151580
rect 180064 29640 180116 29646
rect 180064 29582 180116 29588
rect 175292 16546 175504 16574
rect 176764 16546 177896 16574
rect 178052 16546 178632 16574
rect 179432 16546 180012 16574
rect 174544 3392 174596 3398
rect 174544 3334 174596 3340
rect 175476 480 175504 16546
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 176672 480 176700 3334
rect 177868 480 177896 16546
rect 178040 1692 178092 1698
rect 178040 1634 178092 1640
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178052 66 178080 1634
rect 178604 354 178632 16546
rect 179512 15292 179564 15298
rect 179512 15234 179564 15240
rect 179420 12708 179472 12714
rect 179420 12650 179472 12656
rect 179432 11014 179460 12650
rect 179524 12306 179552 15234
rect 179512 12300 179564 12306
rect 179512 12242 179564 12248
rect 179420 11008 179472 11014
rect 179420 10950 179472 10956
rect 179420 5432 179472 5438
rect 179420 5374 179472 5380
rect 179432 4010 179460 5374
rect 179420 4004 179472 4010
rect 179420 3946 179472 3952
rect 179984 3482 180012 16546
rect 180156 12436 180208 12442
rect 180156 12378 180208 12384
rect 180064 9784 180116 9790
rect 180064 9726 180116 9732
rect 180076 4078 180104 9726
rect 180168 5506 180196 12378
rect 180156 5500 180208 5506
rect 180156 5442 180208 5448
rect 180064 4072 180116 4078
rect 180064 4014 180116 4020
rect 181444 3936 181496 3942
rect 181444 3878 181496 3884
rect 179984 3454 180288 3482
rect 180260 480 180288 3454
rect 181456 480 181484 3878
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 178040 60 178092 66
rect 178040 2 178092 8
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 354 182220 151574
rect 183376 12232 183428 12238
rect 183376 12174 183428 12180
rect 183388 10878 183416 12174
rect 183468 10940 183520 10946
rect 183468 10882 183520 10888
rect 182272 10872 182324 10878
rect 182272 10814 182324 10820
rect 183376 10872 183428 10878
rect 183376 10814 183428 10820
rect 182284 10266 182312 10814
rect 182272 10260 182324 10266
rect 182272 10202 182324 10208
rect 183480 9654 183508 10882
rect 183744 10260 183796 10266
rect 183744 10202 183796 10208
rect 183468 9648 183520 9654
rect 183468 9590 183520 9596
rect 183756 480 183784 10202
rect 184756 8356 184808 8362
rect 184756 8298 184808 8304
rect 184768 6866 184796 8298
rect 184756 6860 184808 6866
rect 184756 6802 184808 6808
rect 184952 3398 184980 154838
rect 188356 24206 188384 162114
rect 196624 162104 196676 162110
rect 196624 162046 196676 162052
rect 191104 158160 191156 158166
rect 191104 158102 191156 158108
rect 191116 156942 191144 158102
rect 191104 156936 191156 156942
rect 191104 156878 191156 156884
rect 192484 156460 192536 156466
rect 192484 156402 192536 156408
rect 189080 151428 189132 151434
rect 189080 151370 189132 151376
rect 188344 24200 188396 24206
rect 188344 24142 188396 24148
rect 187608 18216 187660 18222
rect 187608 18158 187660 18164
rect 187620 15162 187648 18158
rect 189092 16574 189120 151370
rect 192496 150550 192524 156402
rect 192576 156392 192628 156398
rect 192576 156334 192628 156340
rect 192588 151434 192616 156334
rect 195612 154080 195664 154086
rect 195612 154022 195664 154028
rect 195624 151570 195652 154022
rect 193220 151564 193272 151570
rect 193220 151506 193272 151512
rect 195612 151564 195664 151570
rect 195612 151506 195664 151512
rect 192576 151428 192628 151434
rect 192576 151370 192628 151376
rect 192484 150544 192536 150550
rect 192484 150486 192536 150492
rect 190460 24200 190512 24206
rect 190460 24142 190512 24148
rect 189092 16546 189304 16574
rect 187608 15156 187660 15162
rect 187608 15098 187660 15104
rect 188528 14000 188580 14006
rect 188528 13942 188580 13948
rect 186872 8900 186924 8906
rect 186872 8842 186924 8848
rect 186320 6792 186372 6798
rect 186320 6734 186372 6740
rect 185032 5500 185084 5506
rect 185032 5442 185084 5448
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 185044 2802 185072 5442
rect 186332 3942 186360 6734
rect 186884 6118 186912 8842
rect 186872 6112 186924 6118
rect 186872 6054 186924 6060
rect 187332 4072 187384 4078
rect 187332 4014 187384 4020
rect 186320 3936 186372 3942
rect 186320 3878 186372 3884
rect 186136 3392 186188 3398
rect 186136 3334 186188 3340
rect 184952 2774 185072 2802
rect 184952 480 184980 2774
rect 186148 480 186176 3334
rect 187344 480 187372 4014
rect 188540 480 188568 13942
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 24142
rect 191748 8356 191800 8362
rect 191748 8298 191800 8304
rect 191760 7274 191788 8298
rect 191748 7268 191800 7274
rect 191748 7210 191800 7216
rect 191748 6112 191800 6118
rect 191748 6054 191800 6060
rect 191760 3126 191788 6054
rect 192024 4004 192076 4010
rect 192024 3946 192076 3952
rect 191748 3120 191800 3126
rect 191748 3062 191800 3068
rect 192036 480 192064 3946
rect 193232 480 193260 151506
rect 195980 151224 196032 151230
rect 195980 151166 196032 151172
rect 193312 29640 193364 29646
rect 193312 29582 193364 29588
rect 193324 16574 193352 29582
rect 195992 16574 196020 151166
rect 196636 150482 196664 162046
rect 220084 162036 220136 162042
rect 220084 161978 220136 161984
rect 201960 161016 202012 161022
rect 201960 160958 202012 160964
rect 201972 157350 202000 160958
rect 215944 160676 215996 160682
rect 215944 160618 215996 160624
rect 201960 157344 202012 157350
rect 201960 157286 202012 157292
rect 208492 157344 208544 157350
rect 208492 157286 208544 157292
rect 202144 156324 202196 156330
rect 202144 156266 202196 156272
rect 199384 156256 199436 156262
rect 199384 156198 199436 156204
rect 199396 151230 199424 156198
rect 202156 151298 202184 156266
rect 206376 156188 206428 156194
rect 206376 156130 206428 156136
rect 206284 156120 206336 156126
rect 206284 156062 206336 156068
rect 206296 151366 206324 156062
rect 206388 151638 206416 156130
rect 208504 154018 208532 157286
rect 208400 154012 208452 154018
rect 208400 153954 208452 153960
rect 208492 154012 208544 154018
rect 208492 153954 208544 153960
rect 206376 151632 206428 151638
rect 206376 151574 206428 151580
rect 208412 151502 208440 153954
rect 207020 151496 207072 151502
rect 207020 151438 207072 151444
rect 208400 151496 208452 151502
rect 208400 151438 208452 151444
rect 202880 151360 202932 151366
rect 202880 151302 202932 151308
rect 206284 151360 206336 151366
rect 206284 151302 206336 151308
rect 200120 151292 200172 151298
rect 200120 151234 200172 151240
rect 202144 151292 202196 151298
rect 202144 151234 202196 151240
rect 199384 151224 199436 151230
rect 199384 151166 199436 151172
rect 197360 150544 197412 150550
rect 197360 150486 197412 150492
rect 196624 150476 196676 150482
rect 196624 150418 196676 150424
rect 197372 16574 197400 150486
rect 200132 16574 200160 151234
rect 201500 150476 201552 150482
rect 201500 150418 201552 150424
rect 193324 16546 194456 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 200132 16546 200344 16574
rect 194428 480 194456 16546
rect 195980 3868 196032 3874
rect 195980 3810 196032 3816
rect 195612 3120 195664 3126
rect 195612 3062 195664 3068
rect 194968 2984 195020 2990
rect 194968 2926 195020 2932
rect 194980 2174 195008 2926
rect 194968 2168 195020 2174
rect 194968 2110 195020 2116
rect 195624 480 195652 3062
rect 195992 2650 196020 3810
rect 195980 2644 196032 2650
rect 195980 2586 196032 2592
rect 196820 480 196848 16546
rect 197360 14884 197412 14890
rect 197360 14826 197412 14832
rect 197372 12442 197400 14826
rect 197360 12436 197412 12442
rect 197360 12378 197412 12384
rect 197924 480 197952 16546
rect 198740 11008 198792 11014
rect 198740 10950 198792 10956
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 10950
rect 198832 5364 198884 5370
rect 198832 5306 198884 5312
rect 198844 3874 198872 5306
rect 198832 3868 198884 3874
rect 198832 3810 198884 3816
rect 200316 480 200344 16546
rect 201408 16448 201460 16454
rect 201408 16390 201460 16396
rect 201420 13802 201448 16390
rect 201408 13796 201460 13802
rect 201408 13738 201460 13744
rect 200672 3732 200724 3738
rect 200672 3674 200724 3680
rect 200684 2174 200712 3674
rect 201040 2916 201092 2922
rect 201040 2858 201092 2864
rect 200672 2168 200724 2174
rect 200672 2110 200724 2116
rect 201052 2106 201080 2858
rect 201040 2100 201092 2106
rect 201040 2042 201092 2048
rect 201512 480 201540 150418
rect 202892 16574 202920 151302
rect 202892 16546 203472 16574
rect 202696 12436 202748 12442
rect 202696 12378 202748 12384
rect 202236 12164 202288 12170
rect 202236 12106 202288 12112
rect 202248 8158 202276 12106
rect 202236 8152 202288 8158
rect 202236 8094 202288 8100
rect 201684 3800 201736 3806
rect 201684 3742 201736 3748
rect 201696 2106 201724 3742
rect 201684 2100 201736 2106
rect 201684 2042 201736 2048
rect 202708 480 202736 12378
rect 202788 2848 202840 2854
rect 202788 2790 202840 2796
rect 202800 2514 202828 2790
rect 202788 2508 202840 2514
rect 202788 2450 202840 2456
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205088 15156 205140 15162
rect 205088 15098 205140 15104
rect 204168 7948 204220 7954
rect 204168 7890 204220 7896
rect 204180 6118 204208 7890
rect 204812 6860 204864 6866
rect 204812 6802 204864 6808
rect 204168 6112 204220 6118
rect 204168 6054 204220 6060
rect 204824 3738 204852 6802
rect 204812 3732 204864 3738
rect 204812 3674 204864 3680
rect 205100 480 205128 15098
rect 205640 5228 205692 5234
rect 205640 5170 205692 5176
rect 205652 3874 205680 5170
rect 205640 3868 205692 3874
rect 205640 3810 205692 3816
rect 206192 3800 206244 3806
rect 206192 3742 206244 3748
rect 206204 480 206232 3742
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 151438
rect 209778 151328 209834 151337
rect 209778 151263 209834 151272
rect 209792 9674 209820 151263
rect 215956 30326 215984 160618
rect 216036 31068 216088 31074
rect 216036 31010 216088 31016
rect 215944 30320 215996 30326
rect 215944 30262 215996 30268
rect 215300 23996 215352 24002
rect 215300 23938 215352 23944
rect 215312 22778 215340 23938
rect 216048 22846 216076 31010
rect 218060 30320 218112 30326
rect 218060 30262 218112 30268
rect 216036 22840 216088 22846
rect 216036 22782 216088 22788
rect 215300 22772 215352 22778
rect 215300 22714 215352 22720
rect 215300 21276 215352 21282
rect 215300 21218 215352 21224
rect 215312 19990 215340 21218
rect 215300 19984 215352 19990
rect 215300 19926 215352 19932
rect 211068 19848 211120 19854
rect 211068 19790 211120 19796
rect 211080 18630 211108 19790
rect 215300 18828 215352 18834
rect 215300 18770 215352 18776
rect 210056 18624 210108 18630
rect 210056 18566 210108 18572
rect 211068 18624 211120 18630
rect 211068 18566 211120 18572
rect 210068 10946 210096 18566
rect 212816 17672 212868 17678
rect 212816 17614 212868 17620
rect 212828 16454 212856 17614
rect 212816 16448 212868 16454
rect 212816 16390 212868 16396
rect 210976 14952 211028 14958
rect 210976 14894 211028 14900
rect 210988 13054 211016 14894
rect 211804 13728 211856 13734
rect 211804 13670 211856 13676
rect 211068 13660 211120 13666
rect 211068 13602 211120 13608
rect 210976 13048 211028 13054
rect 210976 12990 211028 12996
rect 211080 11490 211108 13602
rect 211068 11484 211120 11490
rect 211068 11426 211120 11432
rect 209872 10940 209924 10946
rect 209872 10882 209924 10888
rect 210056 10940 210108 10946
rect 210056 10882 210108 10888
rect 209700 9646 209820 9674
rect 209700 9586 209728 9646
rect 209688 9580 209740 9586
rect 209688 9522 209740 9528
rect 207664 8084 207716 8090
rect 207664 8026 207716 8032
rect 207676 5234 207704 8026
rect 209884 6914 209912 10882
rect 210976 9580 211028 9586
rect 210976 9522 211028 9528
rect 209792 6886 209912 6914
rect 207664 5228 207716 5234
rect 207664 5170 207716 5176
rect 208584 2848 208636 2854
rect 208584 2790 208636 2796
rect 208596 480 208624 2790
rect 209792 480 209820 6886
rect 210988 480 211016 9522
rect 211816 3806 211844 13670
rect 213368 11484 213420 11490
rect 213368 11426 213420 11432
rect 213000 5296 213052 5302
rect 213000 5238 213052 5244
rect 213012 3942 213040 5238
rect 212172 3936 212224 3942
rect 212172 3878 212224 3884
rect 213000 3936 213052 3942
rect 213000 3878 213052 3884
rect 211804 3800 211856 3806
rect 211804 3742 211856 3748
rect 212184 480 212212 3878
rect 213380 480 213408 11426
rect 213828 8356 213880 8362
rect 213828 8298 213880 8304
rect 213736 8016 213788 8022
rect 213736 7958 213788 7964
rect 213748 6798 213776 7958
rect 213840 7954 213868 8298
rect 213828 7948 213880 7954
rect 213828 7890 213880 7896
rect 213736 6792 213788 6798
rect 213736 6734 213788 6740
rect 214564 6724 214616 6730
rect 214564 6666 214616 6672
rect 214576 5302 214604 6666
rect 214564 5296 214616 5302
rect 214564 5238 214616 5244
rect 214656 3664 214708 3670
rect 214656 3606 214708 3612
rect 214472 2984 214524 2990
rect 214472 2926 214524 2932
rect 214564 2984 214616 2990
rect 214564 2926 214616 2932
rect 214484 480 214512 2926
rect 214576 2718 214604 2926
rect 214668 2718 214696 3606
rect 214564 2712 214616 2718
rect 214564 2654 214616 2660
rect 214656 2712 214708 2718
rect 214656 2654 214708 2660
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 18770
rect 216864 14816 216916 14822
rect 216864 14758 216916 14764
rect 216876 480 216904 14758
rect 218072 11694 218100 30262
rect 220096 28966 220124 161978
rect 233884 161968 233936 161974
rect 233884 161910 233936 161916
rect 233896 30326 233924 161910
rect 285680 161900 285732 161906
rect 285680 161842 285732 161848
rect 246304 160608 246356 160614
rect 246304 160550 246356 160556
rect 238024 157956 238076 157962
rect 238024 157898 238076 157904
rect 238036 30326 238064 157898
rect 233884 30320 233936 30326
rect 233884 30262 233936 30268
rect 236000 30320 236052 30326
rect 236000 30262 236052 30268
rect 238024 30320 238076 30326
rect 238024 30262 238076 30268
rect 240140 30320 240192 30326
rect 240140 30262 240192 30268
rect 220084 28960 220136 28966
rect 220084 28902 220136 28908
rect 222200 28960 222252 28966
rect 222200 28902 222252 28908
rect 218152 22840 218204 22846
rect 218152 22782 218204 22788
rect 218060 11688 218112 11694
rect 218060 11630 218112 11636
rect 218164 6914 218192 22782
rect 222212 16574 222240 28902
rect 222936 19984 222988 19990
rect 222936 19926 222988 19932
rect 222948 19310 222976 19926
rect 222936 19304 222988 19310
rect 222936 19246 222988 19252
rect 226432 19304 226484 19310
rect 226432 19246 226484 19252
rect 222212 16546 222792 16574
rect 222108 12980 222160 12986
rect 222108 12922 222160 12928
rect 222120 12170 222148 12922
rect 222108 12164 222160 12170
rect 222108 12106 222160 12112
rect 219256 11688 219308 11694
rect 219256 11630 219308 11636
rect 218072 6886 218192 6914
rect 218072 480 218100 6886
rect 218152 2848 218204 2854
rect 218152 2790 218204 2796
rect 218164 2446 218192 2790
rect 218152 2440 218204 2446
rect 218152 2382 218204 2388
rect 218244 1488 218296 1494
rect 218244 1430 218296 1436
rect 218256 542 218284 1430
rect 218244 536 218296 542
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 218244 478 218296 484
rect 219268 480 219296 11630
rect 221648 6112 221700 6118
rect 221648 6054 221700 6060
rect 220452 3868 220504 3874
rect 220452 3810 220504 3816
rect 220464 480 220492 3810
rect 221660 3194 221688 6054
rect 221648 3188 221700 3194
rect 221648 3130 221700 3136
rect 220728 3120 220780 3126
rect 220728 3062 220780 3068
rect 220740 2582 220768 3062
rect 221556 2916 221608 2922
rect 221556 2858 221608 2864
rect 220728 2576 220780 2582
rect 220728 2518 220780 2524
rect 221568 480 221596 2858
rect 222764 480 222792 16546
rect 223488 16176 223540 16182
rect 223488 16118 223540 16124
rect 223500 14754 223528 16118
rect 223028 14748 223080 14754
rect 223028 14690 223080 14696
rect 223488 14748 223540 14754
rect 223488 14690 223540 14696
rect 223040 13666 223068 14690
rect 223028 13660 223080 13666
rect 223028 13602 223080 13608
rect 223488 12096 223540 12102
rect 223488 12038 223540 12044
rect 223500 10878 223528 12038
rect 223488 10872 223540 10878
rect 223488 10814 223540 10820
rect 223396 10804 223448 10810
rect 223396 10746 223448 10752
rect 223408 9586 223436 10746
rect 223396 9580 223448 9586
rect 223396 9522 223448 9528
rect 223488 8152 223540 8158
rect 223488 8094 223540 8100
rect 223500 3330 223528 8094
rect 226444 6914 226472 19246
rect 233516 17196 233568 17202
rect 233516 17138 233568 17144
rect 233528 14822 233556 17138
rect 236012 16574 236040 30262
rect 237380 19780 237432 19786
rect 237380 19722 237432 19728
rect 237392 18970 237420 19722
rect 237380 18964 237432 18970
rect 237380 18906 237432 18912
rect 239588 18284 239640 18290
rect 239588 18226 239640 18232
rect 239600 17678 239628 18226
rect 239588 17672 239640 17678
rect 239588 17614 239640 17620
rect 236012 16546 236592 16574
rect 233516 14816 233568 14822
rect 233516 14758 233568 14764
rect 234620 14680 234672 14686
rect 234620 14622 234672 14628
rect 229376 13592 229428 13598
rect 229376 13534 229428 13540
rect 226352 6886 226472 6914
rect 224960 5160 225012 5166
rect 224960 5102 225012 5108
rect 224972 3670 225000 5102
rect 224960 3664 225012 3670
rect 224960 3606 225012 3612
rect 223488 3324 223540 3330
rect 223488 3266 223540 3272
rect 223948 3188 224000 3194
rect 223948 3130 224000 3136
rect 223960 480 223988 3130
rect 225144 2848 225196 2854
rect 225144 2790 225196 2796
rect 225156 480 225184 2790
rect 226352 480 226380 6886
rect 227536 3800 227588 3806
rect 227536 3742 227588 3748
rect 227548 480 227576 3742
rect 228732 1488 228784 1494
rect 228732 1430 228784 1436
rect 228744 480 228772 1430
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 13534
rect 232044 9648 232096 9654
rect 232044 9590 232096 9596
rect 231768 6656 231820 6662
rect 231768 6598 231820 6604
rect 231780 3874 231808 6598
rect 232056 5370 232084 9590
rect 234528 9512 234580 9518
rect 234528 9454 234580 9460
rect 232044 5364 232096 5370
rect 232044 5306 232096 5312
rect 234540 4010 234568 9454
rect 234528 4004 234580 4010
rect 234528 3946 234580 3952
rect 231768 3868 231820 3874
rect 231768 3810 231820 3816
rect 233424 3732 233476 3738
rect 233424 3674 233476 3680
rect 231032 3324 231084 3330
rect 231032 3266 231084 3272
rect 231044 480 231072 3266
rect 232228 3052 232280 3058
rect 232228 2994 232280 3000
rect 232240 480 232268 2994
rect 233436 480 233464 3674
rect 234632 480 234660 14622
rect 236000 10940 236052 10946
rect 236000 10882 236052 10888
rect 236012 9518 236040 10882
rect 236000 9512 236052 9518
rect 236000 9454 236052 9460
rect 236368 7948 236420 7954
rect 236368 7890 236420 7896
rect 236000 5296 236052 5302
rect 236000 5238 236052 5244
rect 236012 3806 236040 5238
rect 236380 5166 236408 7890
rect 236368 5160 236420 5166
rect 236368 5102 236420 5108
rect 236000 3800 236052 3806
rect 236000 3742 236052 3748
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 235828 480 235856 2926
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 238116 3936 238168 3942
rect 238116 3878 238168 3884
rect 237380 2440 237432 2446
rect 237380 2382 237432 2388
rect 237392 610 237420 2382
rect 237380 604 237432 610
rect 237380 546 237432 552
rect 238128 480 238156 3878
rect 239312 1420 239364 1426
rect 239312 1362 239364 1368
rect 239324 480 239352 1362
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 30262
rect 246316 29646 246344 160550
rect 283564 160472 283616 160478
rect 283564 160414 283616 160420
rect 251272 159316 251324 159322
rect 251272 159258 251324 159264
rect 246304 29640 246356 29646
rect 246304 29582 246356 29588
rect 241428 22636 241480 22642
rect 241428 22578 241480 22584
rect 241440 21486 241468 22578
rect 241428 21480 241480 21486
rect 241428 21422 241480 21428
rect 241428 21208 241480 21214
rect 241428 21150 241480 21156
rect 241440 19990 241468 21150
rect 241428 19984 241480 19990
rect 241428 19926 241480 19932
rect 247040 19712 247092 19718
rect 247040 19654 247092 19660
rect 247052 19106 247080 19654
rect 247040 19100 247092 19106
rect 247040 19042 247092 19048
rect 248512 18760 248564 18766
rect 248512 18702 248564 18708
rect 244556 18080 244608 18086
rect 244556 18022 244608 18028
rect 242808 16788 242860 16794
rect 242808 16730 242860 16736
rect 240232 16720 240284 16726
rect 240232 16662 240284 16668
rect 240244 16182 240272 16662
rect 240506 16280 240562 16289
rect 240506 16215 240562 16224
rect 240232 16176 240284 16182
rect 240232 16118 240284 16124
rect 240520 14686 240548 16215
rect 242820 14890 242848 16730
rect 243544 15020 243596 15026
rect 243544 14962 243596 14968
rect 242808 14884 242860 14890
rect 242808 14826 242860 14832
rect 242900 14816 242952 14822
rect 242900 14758 242952 14764
rect 240508 14680 240560 14686
rect 240508 14622 240560 14628
rect 241428 13660 241480 13666
rect 241428 13602 241480 13608
rect 241336 12300 241388 12306
rect 241336 12242 241388 12248
rect 241348 10946 241376 12242
rect 241440 12238 241468 13602
rect 241704 13116 241756 13122
rect 241704 13058 241756 13064
rect 241428 12232 241480 12238
rect 241428 12174 241480 12180
rect 241336 10940 241388 10946
rect 241336 10882 241388 10888
rect 240784 9716 240836 9722
rect 240784 9658 240836 9664
rect 240796 3942 240824 9658
rect 240784 3936 240836 3942
rect 240784 3878 240836 3884
rect 241716 480 241744 13058
rect 242912 3738 242940 14758
rect 243556 13122 243584 14962
rect 244568 14822 244596 18022
rect 244556 14816 244608 14822
rect 244556 14758 244608 14764
rect 244280 13456 244332 13462
rect 244280 13398 244332 13404
rect 243544 13116 243596 13122
rect 243544 13058 243596 13064
rect 244292 12102 244320 13398
rect 244280 12096 244332 12102
rect 244280 12038 244332 12044
rect 248524 11966 248552 18702
rect 251284 16574 251312 159258
rect 267740 159248 267792 159254
rect 267740 159190 267792 159196
rect 253940 29640 253992 29646
rect 253940 29582 253992 29588
rect 253952 16574 253980 29582
rect 255964 26716 256016 26722
rect 255964 26658 256016 26664
rect 254032 23928 254084 23934
rect 254032 23870 254084 23876
rect 254044 19038 254072 23870
rect 255976 22914 256004 26658
rect 255964 22908 256016 22914
rect 255964 22850 256016 22856
rect 260748 21140 260800 21146
rect 260748 21082 260800 21088
rect 254032 19032 254084 19038
rect 254032 18974 254084 18980
rect 260760 18834 260788 21082
rect 266360 19576 266412 19582
rect 266360 19518 266412 19524
rect 266372 19106 266400 19518
rect 260840 19100 260892 19106
rect 260840 19042 260892 19048
rect 266360 19100 266412 19106
rect 266360 19042 266412 19048
rect 260748 18828 260800 18834
rect 260748 18770 260800 18776
rect 260852 16574 260880 19042
rect 263140 18148 263192 18154
rect 263140 18090 263192 18096
rect 251284 16546 251772 16574
rect 253952 16546 254256 16574
rect 260852 16546 261432 16574
rect 249708 12028 249760 12034
rect 249708 11970 249760 11976
rect 245200 11960 245252 11966
rect 245200 11902 245252 11908
rect 248512 11960 248564 11966
rect 248512 11902 248564 11908
rect 242992 9512 243044 9518
rect 242992 9454 243044 9460
rect 242900 3732 242952 3738
rect 242900 3674 242952 3680
rect 243004 3482 243032 9454
rect 244188 3936 244240 3942
rect 244188 3878 244240 3884
rect 244200 3738 244228 3878
rect 244096 3732 244148 3738
rect 244096 3674 244148 3680
rect 244188 3732 244240 3738
rect 244188 3674 244240 3680
rect 242912 3454 243032 3482
rect 242912 480 242940 3454
rect 244108 480 244136 3674
rect 245212 480 245240 11902
rect 249720 10810 249748 11970
rect 249708 10804 249760 10810
rect 249708 10746 249760 10752
rect 249064 10736 249116 10742
rect 249064 10678 249116 10684
rect 247592 5364 247644 5370
rect 247592 5306 247644 5312
rect 246396 3120 246448 3126
rect 246396 3062 246448 3068
rect 246408 480 246436 3062
rect 247040 2848 247092 2854
rect 247040 2790 247092 2796
rect 247052 2446 247080 2790
rect 247040 2440 247092 2446
rect 247040 2382 247092 2388
rect 247604 480 247632 5306
rect 249076 3738 249104 10678
rect 251180 4004 251232 4010
rect 251180 3946 251232 3952
rect 248788 3732 248840 3738
rect 248788 3674 248840 3680
rect 249064 3732 249116 3738
rect 249064 3674 249116 3680
rect 248800 480 248828 3674
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 249996 480 250024 2790
rect 251192 480 251220 3946
rect 251744 3482 251772 16546
rect 253938 16144 253994 16153
rect 253938 16079 253994 16088
rect 251824 14476 251876 14482
rect 251824 14418 251876 14424
rect 251836 4146 251864 14418
rect 253952 13462 253980 16079
rect 253940 13456 253992 13462
rect 253940 13398 253992 13404
rect 251824 4140 251876 4146
rect 251824 4082 251876 4088
rect 252468 4140 252520 4146
rect 252468 4082 252520 4088
rect 251744 3454 252416 3482
rect 252388 480 252416 3454
rect 252480 3330 252508 4082
rect 252468 3324 252520 3330
rect 252468 3266 252520 3272
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 82 253562 480
rect 254228 354 254256 16546
rect 255320 13524 255372 13530
rect 255320 13466 255372 13472
rect 255332 12034 255360 13466
rect 258724 13388 258776 13394
rect 258724 13330 258776 13336
rect 255872 12164 255924 12170
rect 255872 12106 255924 12112
rect 255320 12028 255372 12034
rect 255320 11970 255372 11976
rect 255884 480 255912 12106
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 258276 480 258304 3810
rect 258736 2922 258764 13330
rect 260656 11960 260708 11966
rect 260656 11902 260708 11908
rect 259460 3324 259512 3330
rect 259460 3266 259512 3272
rect 258724 2916 258776 2922
rect 258724 2858 258776 2864
rect 259472 480 259500 3266
rect 260668 480 260696 11902
rect 261404 3482 261432 16546
rect 262496 16380 262548 16386
rect 262496 16322 262548 16328
rect 262508 11966 262536 16322
rect 263152 14482 263180 18090
rect 263600 14884 263652 14890
rect 263600 14826 263652 14832
rect 263140 14476 263192 14482
rect 263140 14418 263192 14424
rect 262496 11960 262548 11966
rect 262496 11902 262548 11908
rect 263612 11898 263640 14826
rect 264980 12028 265032 12034
rect 264980 11970 265032 11976
rect 261484 11892 261536 11898
rect 261484 11834 261536 11840
rect 263600 11892 263652 11898
rect 263600 11834 263652 11840
rect 261496 3874 261524 11834
rect 262864 6180 262916 6186
rect 262864 6122 262916 6128
rect 262876 3942 262904 6122
rect 262864 3936 262916 3942
rect 262864 3878 262916 3884
rect 261484 3868 261536 3874
rect 261484 3810 261536 3816
rect 261404 3454 261800 3482
rect 261772 480 261800 3454
rect 262956 2916 263008 2922
rect 262956 2858 263008 2864
rect 262968 480 262996 2858
rect 264152 2304 264204 2310
rect 264152 2246 264204 2252
rect 264164 480 264192 2246
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 253664 128 253716 134
rect 253450 76 253664 82
rect 253450 70 253716 76
rect 253450 54 253704 70
rect 253450 -960 253562 54
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256700 264 256752 270
rect 257038 218 257150 480
rect 256752 212 257150 218
rect 256700 206 257150 212
rect 256712 190 257150 206
rect 257038 -960 257150 190
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 11970
rect 265624 7880 265676 7886
rect 265624 7822 265676 7828
rect 265636 6186 265664 7822
rect 265624 6180 265676 6186
rect 265624 6122 265676 6128
rect 266544 3868 266596 3874
rect 266544 3810 266596 3816
rect 266556 480 266584 3810
rect 267752 480 267780 159190
rect 278044 149864 278096 149870
rect 278044 149806 278096 149812
rect 278056 41070 278084 149806
rect 278044 41064 278096 41070
rect 278044 41006 278096 41012
rect 282920 41064 282972 41070
rect 282920 41006 282972 41012
rect 282932 36310 282960 41006
rect 283576 40050 283604 160414
rect 283564 40044 283616 40050
rect 283564 39986 283616 39992
rect 282920 36304 282972 36310
rect 282920 36246 282972 36252
rect 284300 22568 284352 22574
rect 284300 22510 284352 22516
rect 284312 21418 284340 22510
rect 284300 21412 284352 21418
rect 284300 21354 284352 21360
rect 270408 19644 270460 19650
rect 270408 19586 270460 19592
rect 267832 18964 267884 18970
rect 267832 18906 267884 18912
rect 267844 16386 267872 18906
rect 270420 18766 270448 19586
rect 276020 19100 276072 19106
rect 276020 19042 276072 19048
rect 270408 18760 270460 18766
rect 270408 18702 270460 18708
rect 270500 18692 270552 18698
rect 270500 18634 270552 18640
rect 270512 16574 270540 18634
rect 270512 16546 270816 16574
rect 267832 16380 267884 16386
rect 267832 16322 267884 16328
rect 270040 12232 270092 12238
rect 270040 12174 270092 12180
rect 268384 10940 268436 10946
rect 268384 10882 268436 10888
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 10882
rect 270052 480 270080 12174
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 276032 13530 276060 19042
rect 280436 19032 280488 19038
rect 280436 18974 280488 18980
rect 280448 16386 280476 18974
rect 283380 18896 283432 18902
rect 283380 18838 283432 18844
rect 280344 16380 280396 16386
rect 280344 16322 280396 16328
rect 280436 16380 280488 16386
rect 280436 16322 280488 16328
rect 276020 13524 276072 13530
rect 276020 13466 276072 13472
rect 280356 13326 280384 16322
rect 283012 16244 283064 16250
rect 283012 16186 283064 16192
rect 282184 14544 282236 14550
rect 282184 14486 282236 14492
rect 282196 13394 282224 14486
rect 282920 13524 282972 13530
rect 282920 13466 282972 13472
rect 282184 13388 282236 13394
rect 282184 13330 282236 13336
rect 276020 13320 276072 13326
rect 276020 13262 276072 13268
rect 280344 13320 280396 13326
rect 280344 13262 280396 13268
rect 276032 10878 276060 13262
rect 276664 10940 276716 10946
rect 276664 10882 276716 10888
rect 276020 10872 276072 10878
rect 276020 10814 276072 10820
rect 272524 6588 272576 6594
rect 272524 6530 272576 6536
rect 272536 3738 272564 6530
rect 274640 5092 274692 5098
rect 274640 5034 274692 5040
rect 273628 3868 273680 3874
rect 273628 3810 273680 3816
rect 272432 3732 272484 3738
rect 272432 3674 272484 3680
rect 272524 3732 272576 3738
rect 272524 3674 272576 3680
rect 272444 480 272472 3674
rect 273640 480 273668 3810
rect 274652 2854 274680 5034
rect 276676 3806 276704 10882
rect 282932 10742 282960 13466
rect 283024 12034 283052 16186
rect 283392 14550 283420 18838
rect 285692 16574 285720 161842
rect 295984 160744 296036 160750
rect 295984 160686 296036 160692
rect 290556 156052 290608 156058
rect 290556 155994 290608 156000
rect 287704 155304 287756 155310
rect 287704 155246 287756 155252
rect 287716 38622 287744 155246
rect 290568 154086 290596 155994
rect 290556 154080 290608 154086
rect 290556 154022 290608 154028
rect 292488 154012 292540 154018
rect 292488 153954 292540 153960
rect 292500 151706 292528 153954
rect 292488 151700 292540 151706
rect 292488 151642 292540 151648
rect 292672 151496 292724 151502
rect 292672 151438 292724 151444
rect 287796 40044 287848 40050
rect 287796 39986 287848 39992
rect 287704 38616 287756 38622
rect 287704 38558 287756 38564
rect 287060 36304 287112 36310
rect 287060 36246 287112 36252
rect 287072 31754 287100 36246
rect 287808 35630 287836 39986
rect 287796 35624 287848 35630
rect 287796 35566 287848 35572
rect 287060 31748 287112 31754
rect 287060 31690 287112 31696
rect 291844 26648 291896 26654
rect 291844 26590 291896 26596
rect 288440 21480 288492 21486
rect 288440 21422 288492 21428
rect 288452 16574 288480 21422
rect 285692 16546 286640 16574
rect 288452 16546 289032 16574
rect 284484 14816 284536 14822
rect 284484 14758 284536 14764
rect 283380 14544 283432 14550
rect 283380 14486 283432 14492
rect 283012 12028 283064 12034
rect 283012 11970 283064 11976
rect 284300 10804 284352 10810
rect 284300 10746 284352 10752
rect 282920 10736 282972 10742
rect 282920 10678 282972 10684
rect 278044 10396 278096 10402
rect 278044 10338 278096 10344
rect 277400 9376 277452 9382
rect 277400 9318 277452 9324
rect 277412 5574 277440 9318
rect 277400 5568 277452 5574
rect 277400 5510 277452 5516
rect 276112 3800 276164 3806
rect 276112 3742 276164 3748
rect 276664 3800 276716 3806
rect 276664 3742 276716 3748
rect 274640 2848 274692 2854
rect 274640 2790 274692 2796
rect 274824 2372 274876 2378
rect 274824 2314 274876 2320
rect 274836 480 274864 2314
rect 276020 1420 276072 1426
rect 276020 1362 276072 1368
rect 276032 746 276060 1362
rect 276020 740 276072 746
rect 276020 682 276072 688
rect 276124 626 276152 3742
rect 277124 3664 277176 3670
rect 277124 3606 277176 3612
rect 276032 598 276152 626
rect 276032 480 276060 598
rect 277136 480 277164 3606
rect 278056 3058 278084 10338
rect 284312 9450 284340 10746
rect 282828 9444 282880 9450
rect 282828 9386 282880 9392
rect 284300 9444 284352 9450
rect 284300 9386 284352 9392
rect 278688 6792 278740 6798
rect 278688 6734 278740 6740
rect 278700 3942 278728 6734
rect 282840 6594 282868 9386
rect 284496 9194 284524 14758
rect 285772 13320 285824 13326
rect 285772 13262 285824 13268
rect 284576 12096 284628 12102
rect 284576 12038 284628 12044
rect 284312 9166 284524 9194
rect 282828 6588 282880 6594
rect 282828 6530 282880 6536
rect 282920 6520 282972 6526
rect 282920 6462 282972 6468
rect 278688 3936 278740 3942
rect 278688 3878 278740 3884
rect 282932 3874 282960 6462
rect 283104 5568 283156 5574
rect 283104 5510 283156 5516
rect 282920 3868 282972 3874
rect 282920 3810 282972 3816
rect 278044 3052 278096 3058
rect 278044 2994 278096 3000
rect 280712 3052 280764 3058
rect 280712 2994 280764 3000
rect 279516 2848 279568 2854
rect 279516 2790 279568 2796
rect 278320 2236 278372 2242
rect 278320 2178 278372 2184
rect 278332 480 278360 2178
rect 279528 480 279556 2790
rect 280724 480 280752 2994
rect 281908 1420 281960 1426
rect 281908 1362 281960 1368
rect 281920 480 281948 1362
rect 283116 480 283144 5510
rect 284312 3670 284340 9166
rect 284588 6914 284616 12038
rect 285680 10668 285732 10674
rect 285680 10610 285732 10616
rect 285692 9382 285720 10610
rect 285784 10402 285812 13262
rect 285772 10396 285824 10402
rect 285772 10338 285824 10344
rect 285680 9376 285732 9382
rect 285680 9318 285732 9324
rect 284404 6886 284616 6914
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 284404 3482 284432 6886
rect 285128 3868 285180 3874
rect 285128 3810 285180 3816
rect 285140 3670 285168 3810
rect 285036 3664 285088 3670
rect 285036 3606 285088 3612
rect 285128 3664 285180 3670
rect 285128 3606 285180 3612
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3606
rect 286612 480 286640 16546
rect 287796 9240 287848 9246
rect 287796 9182 287848 9188
rect 287808 480 287836 9182
rect 289004 480 289032 16546
rect 291752 16312 291804 16318
rect 291752 16254 291804 16260
rect 291764 14890 291792 16254
rect 291752 14884 291804 14890
rect 291752 14826 291804 14832
rect 291752 9308 291804 9314
rect 291752 9250 291804 9256
rect 291764 6526 291792 9250
rect 291752 6520 291804 6526
rect 291752 6462 291804 6468
rect 291752 5024 291804 5030
rect 291752 4966 291804 4972
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 290188 3800 290240 3806
rect 290188 3742 290240 3748
rect 290200 480 290228 3742
rect 291396 480 291424 3810
rect 291764 3806 291792 4966
rect 291752 3800 291804 3806
rect 291752 3742 291804 3748
rect 291856 3126 291884 26590
rect 292212 9580 292264 9586
rect 292212 9522 292264 9528
rect 292224 3874 292252 9522
rect 292684 6914 292712 151438
rect 295340 38616 295392 38622
rect 295340 38558 295392 38564
rect 295352 33794 295380 38558
rect 295996 36582 296024 160686
rect 299492 156874 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 169046 331260 702986
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 331220 169040 331272 169046
rect 331220 168982 331272 168988
rect 302884 161832 302936 161838
rect 302884 161774 302936 161780
rect 300124 159180 300176 159186
rect 300124 159122 300176 159128
rect 299480 156868 299532 156874
rect 299480 156810 299532 156816
rect 295984 36576 296036 36582
rect 295984 36518 296036 36524
rect 295432 35624 295484 35630
rect 295432 35566 295484 35572
rect 295340 33788 295392 33794
rect 295340 33730 295392 33736
rect 295340 31748 295392 31754
rect 295340 31690 295392 31696
rect 295352 28354 295380 31690
rect 295444 29646 295472 35566
rect 300136 35086 300164 159122
rect 300676 36576 300728 36582
rect 300676 36518 300728 36524
rect 300124 35080 300176 35086
rect 300124 35022 300176 35028
rect 299848 33788 299900 33794
rect 299848 33730 299900 33736
rect 295432 29640 295484 29646
rect 295432 29582 295484 29588
rect 299860 28558 299888 33730
rect 300688 32638 300716 36518
rect 302896 33862 302924 161774
rect 305644 161764 305696 161770
rect 305644 161706 305696 161712
rect 303252 35080 303304 35086
rect 303252 35022 303304 35028
rect 302884 33856 302936 33862
rect 302884 33798 302936 33804
rect 300676 32632 300728 32638
rect 300676 32574 300728 32580
rect 302516 32632 302568 32638
rect 302516 32574 302568 32580
rect 299848 28552 299900 28558
rect 299848 28494 299900 28500
rect 302528 28422 302556 32574
rect 303264 31754 303292 35022
rect 305000 33856 305052 33862
rect 305000 33798 305052 33804
rect 303252 31748 303304 31754
rect 303252 31690 303304 31696
rect 305012 29714 305040 33798
rect 305656 32434 305684 161706
rect 309784 161696 309836 161702
rect 309784 161638 309836 161644
rect 305644 32428 305696 32434
rect 305644 32370 305696 32376
rect 309232 32428 309284 32434
rect 309232 32370 309284 32376
rect 305092 31748 305144 31754
rect 305092 31690 305144 31696
rect 305000 29708 305052 29714
rect 305000 29650 305052 29656
rect 305104 28490 305132 31690
rect 305092 28484 305144 28490
rect 305092 28426 305144 28432
rect 302516 28416 302568 28422
rect 302516 28358 302568 28364
rect 295340 28348 295392 28354
rect 295340 28290 295392 28296
rect 309244 28286 309272 32370
rect 309796 31074 309824 161638
rect 353944 160540 353996 160546
rect 353944 160482 353996 160488
rect 336004 160404 336056 160410
rect 336004 160346 336056 160352
rect 331220 157888 331272 157894
rect 331220 157830 331272 157836
rect 323584 156936 323636 156942
rect 323584 156878 323636 156884
rect 317420 154080 317472 154086
rect 317420 154022 317472 154028
rect 317432 151774 317460 154022
rect 323032 152516 323084 152522
rect 323032 152458 323084 152464
rect 317420 151768 317472 151774
rect 317420 151710 317472 151716
rect 319444 151700 319496 151706
rect 319444 151642 319496 151648
rect 313924 149796 313976 149802
rect 313924 149738 313976 149744
rect 309784 31068 309836 31074
rect 309784 31010 309836 31016
rect 309232 28280 309284 28286
rect 309232 28222 309284 28228
rect 303620 25356 303672 25362
rect 303620 25298 303672 25304
rect 303632 24138 303660 25298
rect 303620 24132 303672 24138
rect 303620 24074 303672 24080
rect 305644 23860 305696 23866
rect 305644 23802 305696 23808
rect 300768 21072 300820 21078
rect 300768 21014 300820 21020
rect 300780 20058 300808 21014
rect 300768 20052 300820 20058
rect 300768 19994 300820 20000
rect 299386 19544 299442 19553
rect 299386 19479 299442 19488
rect 299400 18698 299428 19479
rect 302238 18728 302294 18737
rect 299388 18692 299440 18698
rect 302238 18663 302294 18672
rect 299388 18634 299440 18640
rect 294604 17808 294656 17814
rect 294604 17750 294656 17756
rect 294616 16250 294644 17750
rect 302252 16574 302280 18663
rect 302252 16546 303200 16574
rect 295340 16448 295392 16454
rect 295340 16390 295392 16396
rect 294604 16244 294656 16250
rect 294604 16186 294656 16192
rect 295352 14822 295380 16390
rect 298466 14920 298522 14929
rect 298466 14855 298522 14864
rect 295340 14816 295392 14822
rect 295340 14758 295392 14764
rect 297272 14612 297324 14618
rect 297272 14554 297324 14560
rect 292592 6886 292712 6914
rect 292212 3868 292264 3874
rect 292212 3810 292264 3816
rect 291844 3120 291896 3126
rect 291844 3062 291896 3068
rect 292592 480 292620 6886
rect 294972 6452 295024 6458
rect 294972 6394 295024 6400
rect 293684 3732 293736 3738
rect 293684 3674 293736 3680
rect 293696 480 293724 3674
rect 294984 3126 295012 6394
rect 294880 3120 294932 3126
rect 294880 3062 294932 3068
rect 294972 3120 295024 3126
rect 294972 3062 295024 3068
rect 294892 480 294920 3062
rect 297284 480 297312 14554
rect 298480 13326 298508 14855
rect 298468 13320 298520 13326
rect 298468 13262 298520 13268
rect 299388 13048 299440 13054
rect 299388 12990 299440 12996
rect 299400 10674 299428 12990
rect 299480 10872 299532 10878
rect 299480 10814 299532 10820
rect 299388 10668 299440 10674
rect 299388 10610 299440 10616
rect 299492 3398 299520 10814
rect 300768 6384 300820 6390
rect 300768 6326 300820 6332
rect 300780 3738 300808 6326
rect 301964 4956 302016 4962
rect 301964 4898 302016 4904
rect 300768 3732 300820 3738
rect 300768 3674 300820 3680
rect 299480 3392 299532 3398
rect 299480 3334 299532 3340
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 298468 3120 298520 3126
rect 298468 3062 298520 3068
rect 298480 480 298508 3062
rect 299662 2136 299718 2145
rect 299662 2071 299718 2080
rect 299676 480 299704 2071
rect 300780 480 300808 3334
rect 301976 480 302004 4898
rect 303172 480 303200 16546
rect 303620 11824 303672 11830
rect 303620 11766 303672 11772
rect 303632 10810 303660 11766
rect 303620 10804 303672 10810
rect 303620 10746 303672 10752
rect 305552 10600 305604 10606
rect 305552 10542 305604 10548
rect 304356 3664 304408 3670
rect 304356 3606 304408 3612
rect 304368 480 304396 3606
rect 305564 480 305592 10542
rect 305656 3942 305684 23802
rect 309140 23792 309192 23798
rect 309140 23734 309192 23740
rect 306378 18320 306434 18329
rect 306378 18255 306434 18264
rect 305644 3936 305696 3942
rect 305644 3878 305696 3884
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 218 296158 480
rect 295720 202 296158 218
rect 295708 196 296158 202
rect 295760 190 296158 196
rect 295708 138 295760 144
rect 296046 -960 296158 190
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 354 306420 18255
rect 309152 16574 309180 23734
rect 309152 16546 309824 16574
rect 307852 13252 307904 13258
rect 307852 13194 307904 13200
rect 307864 3398 307892 13194
rect 307944 3868 307996 3874
rect 307944 3810 307996 3816
rect 307852 3392 307904 3398
rect 307852 3334 307904 3340
rect 307956 480 307984 3810
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 312176 10804 312228 10810
rect 312176 10746 312228 10752
rect 309876 10668 309928 10674
rect 309876 10610 309928 10616
rect 309888 3874 309916 10610
rect 310428 6316 310480 6322
rect 310428 6258 310480 6264
rect 309876 3868 309928 3874
rect 309876 3810 309928 3816
rect 310440 3670 310468 6258
rect 311440 3800 311492 3806
rect 311440 3742 311492 3748
rect 310428 3664 310480 3670
rect 310428 3606 310480 3612
rect 311452 480 311480 3742
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 10746
rect 313280 10532 313332 10538
rect 313280 10474 313332 10480
rect 313292 9246 313320 10474
rect 313280 9240 313332 9246
rect 313280 9182 313332 9188
rect 313936 4146 313964 149738
rect 318064 26580 318116 26586
rect 318064 26522 318116 26528
rect 317972 14748 318024 14754
rect 317972 14690 318024 14696
rect 314016 13388 314068 13394
rect 314016 13330 314068 13336
rect 314028 5574 314056 13330
rect 317984 6914 318012 14690
rect 318076 13258 318104 26522
rect 318064 13252 318116 13258
rect 318064 13194 318116 13200
rect 318616 13184 318668 13190
rect 318616 13126 318668 13132
rect 318628 7954 318656 13126
rect 318708 9172 318760 9178
rect 318708 9114 318760 9120
rect 318616 7948 318668 7954
rect 318616 7890 318668 7896
rect 318720 7886 318748 9114
rect 318708 7880 318760 7886
rect 318708 7822 318760 7828
rect 317984 6886 318104 6914
rect 314016 5568 314068 5574
rect 314016 5510 314068 5516
rect 316224 5568 316276 5574
rect 316224 5510 316276 5516
rect 315028 5160 315080 5166
rect 315028 5102 315080 5108
rect 313924 4140 313976 4146
rect 313924 4082 313976 4088
rect 313832 3936 313884 3942
rect 313832 3878 313884 3884
rect 313280 1420 313332 1426
rect 313280 1362 313332 1368
rect 313292 1193 313320 1362
rect 313278 1184 313334 1193
rect 313278 1119 313334 1128
rect 313844 480 313872 3878
rect 315040 480 315068 5102
rect 316236 480 316264 5510
rect 317328 4140 317380 4146
rect 317328 4082 317380 4088
rect 317340 480 317368 4082
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 6886
rect 319456 6322 319484 151642
rect 323044 151502 323072 152458
rect 323596 151706 323624 156878
rect 327724 151768 327776 151774
rect 327724 151710 327776 151716
rect 323584 151700 323636 151706
rect 323584 151642 323636 151648
rect 324412 151632 324464 151638
rect 324412 151574 324464 151580
rect 323032 151496 323084 151502
rect 323032 151438 323084 151444
rect 319536 21004 319588 21010
rect 319536 20946 319588 20952
rect 319548 13190 319576 20946
rect 321560 18352 321612 18358
rect 321560 18294 321612 18300
rect 321572 17746 321600 18294
rect 322756 17808 322808 17814
rect 322756 17750 322808 17756
rect 321560 17740 321612 17746
rect 321560 17682 321612 17688
rect 322768 14754 322796 17750
rect 322756 14748 322808 14754
rect 322756 14690 322808 14696
rect 319536 13184 319588 13190
rect 319536 13126 319588 13132
rect 322204 12028 322256 12034
rect 322204 11970 322256 11976
rect 319720 7812 319772 7818
rect 319720 7754 319772 7760
rect 319444 6316 319496 6322
rect 319444 6258 319496 6264
rect 319732 480 319760 7754
rect 321468 7744 321520 7750
rect 321468 7686 321520 7692
rect 321480 3330 321508 7686
rect 321560 6588 321612 6594
rect 321560 6530 321612 6536
rect 321572 3806 321600 6530
rect 321560 3800 321612 3806
rect 321560 3742 321612 3748
rect 322112 3732 322164 3738
rect 322112 3674 322164 3680
rect 321468 3324 321520 3330
rect 321468 3266 321520 3272
rect 320916 1420 320968 1426
rect 320916 1362 320968 1368
rect 320928 480 320956 1362
rect 322124 480 322152 3674
rect 322216 2990 322244 11970
rect 323308 3324 323360 3330
rect 323308 3266 323360 3272
rect 322204 2984 322256 2990
rect 322204 2926 322256 2932
rect 323320 480 323348 3266
rect 324424 480 324452 151574
rect 327736 29782 327764 151710
rect 328092 31068 328144 31074
rect 328092 31010 328144 31016
rect 327724 29776 327776 29782
rect 327724 29718 327776 29724
rect 327816 29708 327868 29714
rect 327816 29650 327868 29656
rect 327080 22500 327132 22506
rect 327080 22442 327132 22448
rect 327092 16574 327120 22442
rect 327828 20126 327856 29650
rect 328104 28626 328132 31010
rect 328092 28620 328144 28626
rect 328092 28562 328144 28568
rect 328000 25288 328052 25294
rect 328000 25230 328052 25236
rect 328012 22846 328040 25230
rect 328000 22840 328052 22846
rect 328000 22782 328052 22788
rect 327816 20120 327868 20126
rect 327816 20062 327868 20068
rect 327092 16546 327672 16574
rect 327540 13796 327592 13802
rect 327540 13738 327592 13744
rect 327552 8294 327580 13738
rect 327540 8288 327592 8294
rect 327540 8230 327592 8236
rect 325608 3868 325660 3874
rect 325608 3810 325660 3816
rect 325620 480 325648 3810
rect 327644 3482 327672 16546
rect 327724 16108 327776 16114
rect 327724 16050 327776 16056
rect 327736 3738 327764 16050
rect 330852 8288 330904 8294
rect 330852 8230 330904 8236
rect 329194 5536 329250 5545
rect 329194 5471 329250 5480
rect 327724 3732 327776 3738
rect 327724 3674 327776 3680
rect 327644 3454 328040 3482
rect 326804 2984 326856 2990
rect 326804 2926 326856 2932
rect 326816 480 326844 2926
rect 328012 480 328040 3454
rect 329208 480 329236 5471
rect 330864 3874 330892 8230
rect 330852 3868 330904 3874
rect 330852 3810 330904 3816
rect 330392 3732 330444 3738
rect 330392 3674 330444 3680
rect 330404 480 330432 3674
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 157830
rect 336016 23322 336044 160346
rect 341524 159044 341576 159050
rect 341524 158986 341576 158992
rect 337384 155236 337436 155242
rect 337384 155178 337436 155184
rect 337396 151638 337424 155178
rect 337384 151632 337436 151638
rect 337384 151574 337436 151580
rect 338120 151564 338172 151570
rect 338120 151506 338172 151512
rect 336096 28620 336148 28626
rect 336096 28562 336148 28568
rect 336004 23316 336056 23322
rect 336004 23258 336056 23264
rect 334624 22908 334676 22914
rect 334624 22850 334676 22856
rect 332692 7948 332744 7954
rect 332692 7890 332744 7896
rect 331312 6316 331364 6322
rect 331312 6258 331364 6264
rect 331324 3806 331352 6258
rect 331312 3800 331364 3806
rect 331312 3742 331364 3748
rect 332704 480 332732 7890
rect 334636 3738 334664 22850
rect 336004 20120 336056 20126
rect 336004 20062 336056 20068
rect 336016 10538 336044 20062
rect 336108 18902 336136 28562
rect 336096 18896 336148 18902
rect 336096 18838 336148 18844
rect 338132 16574 338160 151506
rect 341536 23458 341564 158986
rect 345664 157820 345716 157826
rect 345664 157762 345716 157768
rect 341616 29776 341668 29782
rect 341616 29718 341668 29724
rect 341628 25974 341656 29718
rect 345020 26512 345072 26518
rect 345020 26454 345072 26460
rect 341616 25968 341668 25974
rect 341616 25910 341668 25916
rect 345032 25566 345060 26454
rect 345020 25560 345072 25566
rect 345020 25502 345072 25508
rect 341524 23452 341576 23458
rect 341524 23394 341576 23400
rect 341616 23316 341668 23322
rect 341616 23258 341668 23264
rect 338132 16546 338712 16574
rect 336004 10532 336056 10538
rect 336004 10474 336056 10480
rect 337016 10464 337068 10470
rect 337016 10406 337068 10412
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 334624 3732 334676 3738
rect 334624 3674 334676 3680
rect 333900 480 333928 3674
rect 336280 3664 336332 3670
rect 336280 3606 336332 3612
rect 335082 2000 335138 2009
rect 335082 1935 335138 1944
rect 335096 480 335124 1935
rect 336292 480 336320 3606
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 10406
rect 338684 480 338712 16546
rect 340144 6520 340196 6526
rect 340144 6462 340196 6468
rect 339868 3868 339920 3874
rect 339868 3810 339920 3816
rect 339880 480 339908 3810
rect 340156 3670 340184 6462
rect 341628 6390 341656 23258
rect 345676 22982 345704 157762
rect 349160 157684 349212 157690
rect 349160 157626 349212 157632
rect 346308 25968 346360 25974
rect 346308 25910 346360 25916
rect 345756 23452 345808 23458
rect 345756 23394 345808 23400
rect 345664 22976 345716 22982
rect 345664 22918 345716 22924
rect 343364 9444 343416 9450
rect 343364 9386 343416 9392
rect 342076 7880 342128 7886
rect 342076 7822 342128 7828
rect 341616 6384 341668 6390
rect 341616 6326 341668 6332
rect 340970 5400 341026 5409
rect 340970 5335 341026 5344
rect 340144 3664 340196 3670
rect 340144 3606 340196 3612
rect 340984 480 341012 5335
rect 342088 3874 342116 7822
rect 342076 3868 342128 3874
rect 342076 3810 342128 3816
rect 342168 3800 342220 3806
rect 342168 3742 342220 3748
rect 342180 480 342208 3742
rect 343376 480 343404 9386
rect 345768 6118 345796 23394
rect 346320 22914 346348 25910
rect 346308 22908 346360 22914
rect 346308 22850 346360 22856
rect 345848 22432 345900 22438
rect 345848 22374 345900 22380
rect 345860 7750 345888 22374
rect 349172 16574 349200 157626
rect 350540 149728 350592 149734
rect 350540 149670 350592 149676
rect 349804 28552 349856 28558
rect 349804 28494 349856 28500
rect 349172 16546 349292 16574
rect 348516 11960 348568 11966
rect 348516 11902 348568 11908
rect 348528 9178 348556 11902
rect 348516 9172 348568 9178
rect 348516 9114 348568 9120
rect 345848 7744 345900 7750
rect 345848 7686 345900 7692
rect 345756 6112 345808 6118
rect 345756 6054 345808 6060
rect 346952 5228 347004 5234
rect 346952 5170 347004 5176
rect 344560 3732 344612 3738
rect 344560 3674 344612 3680
rect 344572 480 344600 3674
rect 346964 480 346992 5170
rect 348056 3868 348108 3874
rect 348056 3810 348108 3816
rect 348068 480 348096 3810
rect 349264 480 349292 16546
rect 349816 14958 349844 28494
rect 350552 16574 350580 149670
rect 353956 28558 353984 160482
rect 355324 157752 355376 157758
rect 355324 157694 355376 157700
rect 355336 150482 355364 157694
rect 364352 156806 364380 702406
rect 397472 699718 397500 703520
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 396736 167686 396764 699654
rect 396724 167680 396776 167686
rect 396724 167622 396776 167628
rect 422944 161628 422996 161634
rect 422944 161570 422996 161576
rect 381544 160336 381596 160342
rect 381544 160278 381596 160284
rect 371882 160168 371938 160177
rect 371882 160103 371938 160112
rect 367744 157616 367796 157622
rect 367744 157558 367796 157564
rect 364340 156800 364392 156806
rect 364340 156742 364392 156748
rect 359464 153944 359516 153950
rect 359464 153886 359516 153892
rect 359476 152522 359504 153886
rect 359464 152516 359516 152522
rect 359464 152458 359516 152464
rect 363604 152108 363656 152114
rect 363604 152050 363656 152056
rect 356704 151428 356756 151434
rect 356704 151370 356756 151376
rect 355324 150476 355376 150482
rect 355324 150418 355376 150424
rect 354036 29640 354088 29646
rect 354036 29582 354088 29588
rect 353944 28552 353996 28558
rect 353944 28494 353996 28500
rect 350552 16546 351224 16574
rect 349804 14952 349856 14958
rect 349804 14894 349856 14900
rect 350448 9104 350500 9110
rect 350448 9046 350500 9052
rect 350460 480 350488 9046
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345386 232 345442 241
rect 345726 218 345838 480
rect 345442 190 345838 218
rect 345386 167 345442 176
rect 345726 -960 345838 190
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 353300 14884 353352 14890
rect 353300 14826 353352 14832
rect 351920 13184 351972 13190
rect 351920 13126 351972 13132
rect 351932 8702 351960 13126
rect 353312 11966 353340 14826
rect 353300 11960 353352 11966
rect 353300 11902 353352 11908
rect 354048 10470 354076 29582
rect 355324 26444 355376 26450
rect 355324 26386 355376 26392
rect 355336 13190 355364 26386
rect 355876 25220 355928 25226
rect 355876 25162 355928 25168
rect 355888 21486 355916 25162
rect 355876 21480 355928 21486
rect 355876 21422 355928 21428
rect 355966 16008 356022 16017
rect 355966 15943 356022 15952
rect 355980 14618 356008 15943
rect 355968 14612 356020 14618
rect 355968 14554 356020 14560
rect 355324 13184 355376 13190
rect 355324 13126 355376 13132
rect 354036 10464 354088 10470
rect 354036 10406 354088 10412
rect 356716 9586 356744 151370
rect 359464 150476 359516 150482
rect 359464 150418 359516 150424
rect 359476 23050 359504 150418
rect 359556 28484 359608 28490
rect 359556 28426 359608 28432
rect 359464 23044 359516 23050
rect 359464 22986 359516 22992
rect 356796 22976 356848 22982
rect 356796 22918 356848 22924
rect 356808 9654 356836 22918
rect 358726 14784 358782 14793
rect 358726 14719 358782 14728
rect 358740 12034 358768 14719
rect 358728 12028 358780 12034
rect 358728 11970 358780 11976
rect 356796 9648 356848 9654
rect 356796 9590 356848 9596
rect 356704 9580 356756 9586
rect 356704 9522 356756 9528
rect 354036 9376 354088 9382
rect 354036 9318 354088 9324
rect 351920 8696 351972 8702
rect 351920 8638 351972 8644
rect 353022 8256 353078 8265
rect 353022 8191 353078 8200
rect 353036 6322 353064 8191
rect 353024 6316 353076 6322
rect 353024 6258 353076 6264
rect 351920 6112 351972 6118
rect 351920 6054 351972 6060
rect 351932 3670 351960 6054
rect 352840 3732 352892 3738
rect 352840 3674 352892 3680
rect 351920 3664 351972 3670
rect 351920 3606 351972 3612
rect 352852 480 352880 3674
rect 354048 480 354076 9318
rect 357532 9172 357584 9178
rect 357532 9114 357584 9120
rect 355232 9036 355284 9042
rect 355232 8978 355284 8984
rect 354680 8696 354732 8702
rect 354680 8638 354732 8644
rect 354692 3398 354720 8638
rect 354680 3392 354732 3398
rect 354680 3334 354732 3340
rect 355244 480 355272 8978
rect 357544 480 357572 9114
rect 358818 6760 358874 6769
rect 358818 6695 358874 6704
rect 358832 3398 358860 6695
rect 359568 6458 359596 28426
rect 363616 13394 363644 152050
rect 363696 23044 363748 23050
rect 363696 22986 363748 22992
rect 363604 13388 363656 13394
rect 363604 13330 363656 13336
rect 362960 10532 363012 10538
rect 362960 10474 363012 10480
rect 360108 9648 360160 9654
rect 360108 9590 360160 9596
rect 360016 9580 360068 9586
rect 360016 9522 360068 9528
rect 359556 6452 359608 6458
rect 359556 6394 359608 6400
rect 360028 6118 360056 9522
rect 360016 6112 360068 6118
rect 360016 6054 360068 6060
rect 359924 3664 359976 3670
rect 359924 3606 359976 3612
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358820 3392 358872 3398
rect 358820 3334 358872 3340
rect 358740 480 358768 3334
rect 359936 480 359964 3606
rect 360120 3194 360148 9590
rect 362972 7818 363000 10474
rect 362960 7812 363012 7818
rect 362960 7754 363012 7760
rect 363052 6384 363104 6390
rect 363052 6326 363104 6332
rect 361120 6248 361172 6254
rect 361120 6190 361172 6196
rect 360108 3188 360160 3194
rect 360108 3130 360160 3136
rect 361132 480 361160 6190
rect 362960 6112 363012 6118
rect 362960 6054 363012 6060
rect 362972 4146 363000 6054
rect 362960 4140 363012 4146
rect 362960 4082 363012 4088
rect 362316 3392 362368 3398
rect 362316 3334 362368 3340
rect 362328 480 362356 3334
rect 363064 2922 363092 6326
rect 363708 6254 363736 22986
rect 367650 14648 367706 14657
rect 367650 14583 367706 14592
rect 364616 7676 364668 7682
rect 364616 7618 364668 7624
rect 363696 6248 363748 6254
rect 363696 6190 363748 6196
rect 363512 3188 363564 3194
rect 363512 3130 363564 3136
rect 363052 2916 363104 2922
rect 363052 2858 363104 2864
rect 363524 480 363552 3130
rect 364628 480 364656 7618
rect 367664 6914 367692 14583
rect 367756 9654 367784 157558
rect 368480 155984 368532 155990
rect 368480 155926 368532 155932
rect 368492 16574 368520 155926
rect 371896 35894 371924 160103
rect 374000 158976 374052 158982
rect 374000 158918 374052 158924
rect 371896 35866 372016 35894
rect 371884 28348 371936 28354
rect 371884 28290 371936 28296
rect 371896 25634 371924 28290
rect 371884 25628 371936 25634
rect 371884 25570 371936 25576
rect 371988 22982 372016 35866
rect 371976 22976 372028 22982
rect 371976 22918 372028 22924
rect 371240 22908 371292 22914
rect 371240 22850 371292 22856
rect 370504 21480 370556 21486
rect 370504 21422 370556 21428
rect 368492 16546 369440 16574
rect 367836 10464 367888 10470
rect 367836 10406 367888 10412
rect 367744 9648 367796 9654
rect 367744 9590 367796 9596
rect 367664 6886 367784 6914
rect 367008 4140 367060 4146
rect 367008 4082 367060 4088
rect 365812 2916 365864 2922
rect 365812 2858 365864 2864
rect 365824 480 365852 2858
rect 367020 480 367048 4082
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 82 356418 480
rect 356306 66 356560 82
rect 356306 60 356572 66
rect 356306 54 356520 60
rect 356306 -960 356418 54
rect 356520 2 356572 8
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 6886
rect 367848 5710 367876 10406
rect 368388 6248 368440 6254
rect 368388 6190 368440 6196
rect 367836 5704 367888 5710
rect 367836 5646 367888 5652
rect 368400 2922 368428 6190
rect 368388 2916 368440 2922
rect 368388 2858 368440 2864
rect 369412 480 369440 16546
rect 370516 6254 370544 21422
rect 371252 20126 371280 22850
rect 371240 20120 371292 20126
rect 371240 20062 371292 20068
rect 373264 17740 373316 17746
rect 373264 17682 373316 17688
rect 372620 17604 372672 17610
rect 372620 17546 372672 17552
rect 372632 16114 372660 17546
rect 372620 16108 372672 16114
rect 372620 16050 372672 16056
rect 371238 13288 371294 13297
rect 371238 13223 371294 13232
rect 370504 6248 370556 6254
rect 370504 6190 370556 6196
rect 370964 5704 371016 5710
rect 370964 5646 371016 5652
rect 370976 3738 371004 5646
rect 370964 3732 371016 3738
rect 370964 3674 371016 3680
rect 370596 2916 370648 2922
rect 370596 2858 370648 2864
rect 370608 480 370636 2858
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 13223
rect 372896 9648 372948 9654
rect 372896 9590 372948 9596
rect 372618 6624 372674 6633
rect 372618 6559 372674 6568
rect 372632 3330 372660 6559
rect 372620 3324 372672 3330
rect 372620 3266 372672 3272
rect 372908 480 372936 9590
rect 373276 6390 373304 17682
rect 373264 6384 373316 6390
rect 373264 6326 373316 6332
rect 374012 1170 374040 158918
rect 377404 151700 377456 151706
rect 377404 151642 377456 151648
rect 377416 19310 377444 151642
rect 377956 28416 378008 28422
rect 377956 28358 378008 28364
rect 377968 22914 377996 28358
rect 380900 25628 380952 25634
rect 380900 25570 380952 25576
rect 378048 22976 378100 22982
rect 378048 22918 378100 22924
rect 377956 22908 378008 22914
rect 377956 22850 378008 22856
rect 378060 20126 378088 22918
rect 380912 20194 380940 25570
rect 381556 24206 381584 160278
rect 400220 160268 400272 160274
rect 400220 160210 400272 160216
rect 386420 159112 386472 159118
rect 386420 159054 386472 159060
rect 385684 158840 385736 158846
rect 385684 158782 385736 158788
rect 385696 30326 385724 158782
rect 385684 30320 385736 30326
rect 385684 30262 385736 30268
rect 381636 28552 381688 28558
rect 381636 28494 381688 28500
rect 381544 24200 381596 24206
rect 381544 24142 381596 24148
rect 380900 20188 380952 20194
rect 380900 20130 380952 20136
rect 377588 20120 377640 20126
rect 377588 20062 377640 20068
rect 378048 20120 378100 20126
rect 378048 20062 378100 20068
rect 377404 19304 377456 19310
rect 377404 19246 377456 19252
rect 374092 16040 374144 16046
rect 374092 15982 374144 15988
rect 374104 3398 374132 15982
rect 377600 15366 377628 20062
rect 381544 18896 381596 18902
rect 381544 18838 381596 18844
rect 378048 17536 378100 17542
rect 378048 17478 378100 17484
rect 377772 16108 377824 16114
rect 377772 16050 377824 16056
rect 377588 15360 377640 15366
rect 377588 15302 377640 15308
rect 377784 12442 377812 16050
rect 377772 12436 377824 12442
rect 377772 12378 377824 12384
rect 378060 12170 378088 17478
rect 380900 16380 380952 16386
rect 380900 16322 380952 16328
rect 378048 12164 378100 12170
rect 378048 12106 378100 12112
rect 377954 11928 378010 11937
rect 377954 11863 378010 11872
rect 377402 10568 377458 10577
rect 377402 10503 377458 10512
rect 377416 3670 377444 10503
rect 377680 9240 377732 9246
rect 377680 9182 377732 9188
rect 377404 3664 377456 3670
rect 377404 3606 377456 3612
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 376484 3324 376536 3330
rect 376484 3266 376536 3272
rect 376496 480 376524 3266
rect 377692 480 377720 9182
rect 377968 9042 377996 11863
rect 380912 11830 380940 16322
rect 381556 16114 381584 18838
rect 381648 17542 381676 28494
rect 381912 19304 381964 19310
rect 381912 19246 381964 19252
rect 381636 17536 381688 17542
rect 381636 17478 381688 17484
rect 381544 16108 381596 16114
rect 381544 16050 381596 16056
rect 381924 16046 381952 19246
rect 386432 16574 386460 159054
rect 388444 158908 388496 158914
rect 388444 158850 388496 158856
rect 388456 28354 388484 158850
rect 391204 157548 391256 157554
rect 391204 157490 391256 157496
rect 388536 30320 388588 30326
rect 388536 30262 388588 30268
rect 388444 28348 388496 28354
rect 388444 28290 388496 28296
rect 388548 24682 388576 30262
rect 388536 24676 388588 24682
rect 388536 24618 388588 24624
rect 388352 24200 388404 24206
rect 388352 24142 388404 24148
rect 388364 18902 388392 24142
rect 391216 22914 391244 157490
rect 394700 151360 394752 151366
rect 394700 151302 394752 151308
rect 391296 24676 391348 24682
rect 391296 24618 391348 24624
rect 388536 22908 388588 22914
rect 388536 22850 388588 22856
rect 391204 22908 391256 22914
rect 391204 22850 391256 22856
rect 388352 18896 388404 18902
rect 388352 18838 388404 18844
rect 388444 18828 388496 18834
rect 388444 18770 388496 18776
rect 386432 16546 386736 16574
rect 381912 16040 381964 16046
rect 381912 15982 381964 15988
rect 381176 15360 381228 15366
rect 381176 15302 381228 15308
rect 380992 12436 381044 12442
rect 380992 12378 381044 12384
rect 380900 11824 380952 11830
rect 380900 11766 380952 11772
rect 378048 11212 378100 11218
rect 378048 11154 378100 11160
rect 378060 9110 378088 11154
rect 381004 9178 381032 12378
rect 380992 9172 381044 9178
rect 380992 9114 381044 9120
rect 378048 9104 378100 9110
rect 378048 9046 378100 9052
rect 377956 9036 378008 9042
rect 377956 8978 378008 8984
rect 378874 6488 378930 6497
rect 378874 6423 378930 6432
rect 378888 480 378916 6423
rect 379980 3732 380032 3738
rect 379980 3674 380032 3680
rect 379992 480 380020 3674
rect 381188 480 381216 15302
rect 385314 10432 385370 10441
rect 385314 10367 385370 10376
rect 385328 8974 385356 10367
rect 382372 8968 382424 8974
rect 382372 8910 382424 8916
rect 385316 8968 385368 8974
rect 385316 8910 385368 8916
rect 382384 480 382412 8910
rect 383568 7744 383620 7750
rect 383568 7686 383620 7692
rect 383580 480 383608 7686
rect 385960 7608 386012 7614
rect 385960 7550 386012 7556
rect 384394 912 384450 921
rect 384394 847 384450 856
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384408 354 384436 847
rect 385972 480 386000 7550
rect 384734 354 384846 480
rect 384408 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387800 11824 387852 11830
rect 387800 11766 387852 11772
rect 387812 9654 387840 11766
rect 387800 9648 387852 9654
rect 387800 9590 387852 9596
rect 388456 3670 388484 18770
rect 388548 12442 388576 22850
rect 391308 16318 391336 24618
rect 394712 16574 394740 151302
rect 399484 151292 399536 151298
rect 399484 151234 399536 151240
rect 395344 28280 395396 28286
rect 395344 28222 395396 28228
rect 394712 16546 395292 16574
rect 391296 16312 391348 16318
rect 391296 16254 391348 16260
rect 390652 16040 390704 16046
rect 390652 15982 390704 15988
rect 390560 14952 390612 14958
rect 390560 14894 390612 14900
rect 388536 12436 388588 12442
rect 388536 12378 388588 12384
rect 390572 11830 390600 14894
rect 390560 11824 390612 11830
rect 390560 11766 390612 11772
rect 389088 7812 389140 7818
rect 389088 7754 389140 7760
rect 389100 3738 389128 7754
rect 390664 6914 390692 15982
rect 390928 12436 390980 12442
rect 390928 12378 390980 12384
rect 390940 9246 390968 12378
rect 394976 12164 395028 12170
rect 394976 12106 395028 12112
rect 391848 9648 391900 9654
rect 391848 9590 391900 9596
rect 390928 9240 390980 9246
rect 390928 9182 390980 9188
rect 390572 6886 390692 6914
rect 389454 5264 389510 5273
rect 389454 5199 389510 5208
rect 389088 3732 389140 3738
rect 389088 3674 389140 3680
rect 388260 3664 388312 3670
rect 388260 3606 388312 3612
rect 388444 3664 388496 3670
rect 388444 3606 388496 3612
rect 388272 480 388300 3606
rect 389468 480 389496 5199
rect 390572 3398 390600 6886
rect 391860 6730 391888 9590
rect 394988 9110 395016 12106
rect 393044 9104 393096 9110
rect 393044 9046 393096 9052
rect 394976 9104 395028 9110
rect 394976 9046 395028 9052
rect 391848 6724 391900 6730
rect 391848 6666 391900 6672
rect 390652 6452 390704 6458
rect 390652 6394 390704 6400
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 6394
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 393056 480 393084 9046
rect 394700 8968 394752 8974
rect 394700 8910 394752 8916
rect 394712 5574 394740 8910
rect 395264 6914 395292 16546
rect 395356 16046 395384 28222
rect 399496 23458 399524 151234
rect 400036 28348 400088 28354
rect 400036 28290 400088 28296
rect 399484 23452 399536 23458
rect 399484 23394 399536 23400
rect 399576 22364 399628 22370
rect 399576 22306 399628 22312
rect 399484 20188 399536 20194
rect 399484 20130 399536 20136
rect 399024 16312 399076 16318
rect 399024 16254 399076 16260
rect 395804 16108 395856 16114
rect 395804 16050 395856 16056
rect 395344 16040 395396 16046
rect 395344 15982 395396 15988
rect 395816 12102 395844 16050
rect 396080 14680 396132 14686
rect 396080 14622 396132 14628
rect 395804 12096 395856 12102
rect 395804 12038 395856 12044
rect 395264 6886 395384 6914
rect 394700 5568 394752 5574
rect 394700 5510 394752 5516
rect 394240 3732 394292 3738
rect 394240 3674 394292 3680
rect 394252 480 394280 3674
rect 395356 480 395384 6886
rect 395436 6724 395488 6730
rect 395436 6666 395488 6672
rect 395448 3058 395476 6666
rect 395436 3052 395488 3058
rect 395436 2994 395488 3000
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 14622
rect 398932 13388 398984 13394
rect 398932 13330 398984 13336
rect 398840 11144 398892 11150
rect 398840 11086 398892 11092
rect 398852 8974 398880 11086
rect 398944 10538 398972 13330
rect 398932 10532 398984 10538
rect 398932 10474 398984 10480
rect 398840 8968 398892 8974
rect 398840 8910 398892 8916
rect 399036 6914 399064 16254
rect 399496 16114 399524 20130
rect 399484 16108 399536 16114
rect 399484 16050 399536 16056
rect 399588 14890 399616 22306
rect 400048 20194 400076 28290
rect 400036 20188 400088 20194
rect 400036 20130 400088 20136
rect 400232 16574 400260 160210
rect 421564 158772 421616 158778
rect 421564 158714 421616 158720
rect 417424 157480 417476 157486
rect 417424 157422 417476 157428
rect 409144 153876 409196 153882
rect 409144 153818 409196 153824
rect 406384 152516 406436 152522
rect 406384 152458 406436 152464
rect 403624 151632 403676 151638
rect 403624 151574 403676 151580
rect 403636 23798 403664 151574
rect 406396 27606 406424 152458
rect 406384 27600 406436 27606
rect 406384 27542 406436 27548
rect 409052 27600 409104 27606
rect 409052 27542 409104 27548
rect 403900 25152 403952 25158
rect 403900 25094 403952 25100
rect 403624 23792 403676 23798
rect 403624 23734 403676 23740
rect 403624 23452 403676 23458
rect 403624 23394 403676 23400
rect 400232 16546 400904 16574
rect 399576 14884 399628 14890
rect 399576 14826 399628 14832
rect 400128 9240 400180 9246
rect 400128 9182 400180 9188
rect 398944 6886 399064 6914
rect 397736 3052 397788 3058
rect 397736 2994 397788 3000
rect 397748 480 397776 2994
rect 398944 480 398972 6886
rect 400140 6594 400168 9182
rect 400128 6588 400180 6594
rect 400128 6530 400180 6536
rect 400128 5568 400180 5574
rect 400128 5510 400180 5516
rect 400140 480 400168 5510
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 403636 9654 403664 23394
rect 403716 20120 403768 20126
rect 403716 20062 403768 20068
rect 403728 12442 403756 20062
rect 403912 18834 403940 25094
rect 406660 23792 406712 23798
rect 406660 23734 406712 23740
rect 406672 20670 406700 23734
rect 409064 23050 409092 27542
rect 409156 26110 409184 153818
rect 409144 26104 409196 26110
rect 409144 26046 409196 26052
rect 413468 26104 413520 26110
rect 413468 26046 413520 26052
rect 409052 23044 409104 23050
rect 409052 22986 409104 22992
rect 408592 22908 408644 22914
rect 408592 22850 408644 22856
rect 406660 20664 406712 20670
rect 406660 20606 406712 20612
rect 407028 20188 407080 20194
rect 407028 20130 407080 20136
rect 403900 18828 403952 18834
rect 403900 18770 403952 18776
rect 407040 17610 407068 20130
rect 408604 18766 408632 22850
rect 413480 22370 413508 26046
rect 417436 22914 417464 157422
rect 421576 23050 421604 158714
rect 422956 151298 422984 161570
rect 429212 156738 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 164898 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 462320 164892 462372 164898
rect 462320 164834 462372 164840
rect 449164 161560 449216 161566
rect 449164 161502 449216 161508
rect 445024 160200 445076 160206
rect 445024 160142 445076 160148
rect 429200 156732 429252 156738
rect 429200 156674 429252 156680
rect 427084 155712 427136 155718
rect 427084 155654 427136 155660
rect 427096 153882 427124 155654
rect 442262 155136 442318 155145
rect 442262 155071 442318 155080
rect 439502 154184 439558 154193
rect 439502 154119 439558 154128
rect 427084 153876 427136 153882
rect 427084 153818 427136 153824
rect 427084 153604 427136 153610
rect 427084 153546 427136 153552
rect 422944 151292 422996 151298
rect 422944 151234 422996 151240
rect 417516 23044 417568 23050
rect 417516 22986 417568 22992
rect 421564 23044 421616 23050
rect 421564 22986 421616 22992
rect 426808 23044 426860 23050
rect 426808 22986 426860 22992
rect 417424 22908 417476 22914
rect 417424 22850 417476 22856
rect 413468 22364 413520 22370
rect 413468 22306 413520 22312
rect 413928 20936 413980 20942
rect 413928 20878 413980 20884
rect 413284 20664 413336 20670
rect 413284 20606 413336 20612
rect 408500 18760 408552 18766
rect 408500 18702 408552 18708
rect 408592 18760 408644 18766
rect 408592 18702 408644 18708
rect 407028 17604 407080 17610
rect 407028 17546 407080 17552
rect 406566 17368 406622 17377
rect 406566 17303 406622 17312
rect 406580 14686 406608 17303
rect 408512 16574 408540 18702
rect 412640 17468 412692 17474
rect 412640 17410 412692 17416
rect 408512 16546 409184 16574
rect 407120 14816 407172 14822
rect 407120 14758 407172 14764
rect 406568 14680 406620 14686
rect 406568 14622 406620 14628
rect 405832 13320 405884 13326
rect 405832 13262 405884 13268
rect 403716 12436 403768 12442
rect 403716 12378 403768 12384
rect 404266 11792 404322 11801
rect 404266 11727 404322 11736
rect 403624 9648 403676 9654
rect 403624 9590 403676 9596
rect 403714 9344 403770 9353
rect 404280 9314 404308 11727
rect 405844 9586 405872 13262
rect 406016 9648 406068 9654
rect 406016 9590 406068 9596
rect 405832 9580 405884 9586
rect 405832 9522 405884 9528
rect 403714 9279 403770 9288
rect 404268 9308 404320 9314
rect 403164 9104 403216 9110
rect 403164 9046 403216 9052
rect 403176 6322 403204 9046
rect 403532 6384 403584 6390
rect 403532 6326 403584 6332
rect 403164 6316 403216 6322
rect 403164 6258 403216 6264
rect 402520 3664 402572 3670
rect 402520 3606 402572 3612
rect 402532 480 402560 3606
rect 403544 3210 403572 6326
rect 403728 6254 403756 9279
rect 404268 9250 404320 9256
rect 403624 6248 403676 6254
rect 403624 6190 403676 6196
rect 403716 6248 403768 6254
rect 403716 6190 403768 6196
rect 403636 3670 403664 6190
rect 403624 3664 403676 3670
rect 403624 3606 403676 3612
rect 403544 3182 403664 3210
rect 403636 480 403664 3182
rect 404820 2168 404872 2174
rect 404820 2110 404872 2116
rect 404832 480 404860 2110
rect 406028 480 406056 9590
rect 407132 3398 407160 14758
rect 408500 12436 408552 12442
rect 408500 12378 408552 12384
rect 408512 9246 408540 12378
rect 408684 9580 408736 9586
rect 408684 9522 408736 9528
rect 408500 9240 408552 9246
rect 408500 9182 408552 9188
rect 408696 6458 408724 9522
rect 408684 6452 408736 6458
rect 408684 6394 408736 6400
rect 407210 6352 407266 6361
rect 407210 6287 407266 6296
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 6287
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410798 15872 410854 15881
rect 410798 15807 410854 15816
rect 409788 2848 409840 2854
rect 409788 2790 409840 2796
rect 409800 2650 409828 2790
rect 409788 2644 409840 2650
rect 409788 2586 409840 2592
rect 410812 480 410840 15807
rect 412652 14822 412680 17410
rect 412640 14816 412692 14822
rect 412640 14758 412692 14764
rect 412640 9172 412692 9178
rect 412640 9114 412692 9120
rect 412652 5574 412680 9114
rect 413100 6520 413152 6526
rect 413100 6462 413152 6468
rect 412640 5568 412692 5574
rect 412640 5510 412692 5516
rect 411904 2848 411956 2854
rect 411904 2790 411956 2796
rect 411916 480 411944 2790
rect 413112 480 413140 6462
rect 413296 3194 413324 20606
rect 413940 20126 413968 20878
rect 413928 20120 413980 20126
rect 413928 20062 413980 20068
rect 417424 18760 417476 18766
rect 417424 18702 417476 18708
rect 417332 16244 417384 16250
rect 417332 16186 417384 16192
rect 413560 14884 413612 14890
rect 413560 14826 413612 14832
rect 413572 9110 413600 14826
rect 417240 13184 417292 13190
rect 417240 13126 417292 13132
rect 417252 10470 417280 13126
rect 417344 12238 417372 16186
rect 417436 14142 417464 18702
rect 417528 17066 417556 22986
rect 421012 22364 421064 22370
rect 421012 22306 421064 22312
rect 421024 17610 421052 22306
rect 424968 21412 425020 21418
rect 424968 21354 425020 21360
rect 424980 17950 425008 21354
rect 424968 17944 425020 17950
rect 424968 17886 425020 17892
rect 420920 17604 420972 17610
rect 420920 17546 420972 17552
rect 421012 17604 421064 17610
rect 421012 17546 421064 17552
rect 417516 17060 417568 17066
rect 417516 17002 417568 17008
rect 420932 14210 420960 17546
rect 426820 17406 426848 22986
rect 422392 17400 422444 17406
rect 422392 17342 422444 17348
rect 426808 17400 426860 17406
rect 426808 17342 426860 17348
rect 422404 16574 422432 17342
rect 423680 17060 423732 17066
rect 423680 17002 423732 17008
rect 422404 16546 422616 16574
rect 420920 14204 420972 14210
rect 420920 14146 420972 14152
rect 417424 14136 417476 14142
rect 417424 14078 417476 14084
rect 420918 13152 420974 13161
rect 420918 13087 420974 13096
rect 417332 12232 417384 12238
rect 417332 12174 417384 12180
rect 417424 10736 417476 10742
rect 417424 10678 417476 10684
rect 417240 10464 417292 10470
rect 417240 10406 417292 10412
rect 414294 9208 414350 9217
rect 414294 9143 414350 9152
rect 413560 9104 413612 9110
rect 413560 9046 413612 9052
rect 413284 3188 413336 3194
rect 413284 3130 413336 3136
rect 414308 480 414336 9143
rect 416872 8968 416924 8974
rect 416872 8910 416924 8916
rect 416884 6390 416912 8910
rect 417436 6526 417464 10678
rect 417424 6520 417476 6526
rect 417424 6462 417476 6468
rect 417884 6452 417936 6458
rect 417884 6394 417936 6400
rect 416872 6384 416924 6390
rect 416872 6326 416924 6332
rect 415492 5568 415544 5574
rect 415492 5510 415544 5516
rect 415504 480 415532 5510
rect 416688 3188 416740 3194
rect 416688 3130 416740 3136
rect 416700 480 416728 3130
rect 417896 480 417924 6394
rect 420184 3664 420236 3670
rect 420184 3606 420236 3612
rect 418988 2100 419040 2106
rect 418988 2042 419040 2048
rect 419000 480 419028 2042
rect 420196 480 420224 3606
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 13087
rect 421564 11892 421616 11898
rect 421564 11834 421616 11840
rect 421576 6458 421604 11834
rect 421564 6452 421616 6458
rect 421564 6394 421616 6400
rect 422588 480 422616 16546
rect 423692 14822 423720 17002
rect 427096 16574 427124 153546
rect 431224 153536 431276 153542
rect 431224 153478 431276 153484
rect 430580 22908 430632 22914
rect 430580 22850 430632 22856
rect 430592 20194 430620 22850
rect 430580 20188 430632 20194
rect 430580 20130 430632 20136
rect 431236 17610 431264 153478
rect 435364 151292 435416 151298
rect 435364 151234 435416 151240
rect 431316 17944 431368 17950
rect 431316 17886 431368 17892
rect 427636 17604 427688 17610
rect 427636 17546 427688 17552
rect 431224 17604 431276 17610
rect 431224 17546 431276 17552
rect 427004 16546 427124 16574
rect 423588 14816 423640 14822
rect 423588 14758 423640 14764
rect 423680 14816 423732 14822
rect 423680 14758 423732 14764
rect 423600 12374 423628 14758
rect 424968 14204 425020 14210
rect 424968 14146 425020 14152
rect 423772 14136 423824 14142
rect 423772 14078 423824 14084
rect 423588 12368 423640 12374
rect 423588 12310 423640 12316
rect 423784 480 423812 14078
rect 424980 9178 425008 14146
rect 424968 9172 425020 9178
rect 424968 9114 425020 9120
rect 427004 8974 427032 16546
rect 427648 14686 427676 17546
rect 427084 14680 427136 14686
rect 427084 14622 427136 14628
rect 427636 14680 427688 14686
rect 427636 14622 427688 14628
rect 427096 12170 427124 14622
rect 430578 14512 430634 14521
rect 430578 14447 430634 14456
rect 430592 12306 430620 14447
rect 430580 12300 430632 12306
rect 430580 12242 430632 12248
rect 427084 12164 427136 12170
rect 427084 12106 427136 12112
rect 427176 10532 427228 10538
rect 427176 10474 427228 10480
rect 426992 8968 427044 8974
rect 426992 8910 427044 8916
rect 424966 8120 425022 8129
rect 424966 8055 425022 8064
rect 424980 480 425008 8055
rect 427188 6390 427216 10474
rect 427728 9308 427780 9314
rect 427728 9250 427780 9256
rect 427740 6662 427768 9250
rect 431328 9042 431356 17886
rect 435376 17474 435404 151234
rect 438860 22296 438912 22302
rect 438860 22238 438912 22244
rect 435548 20188 435600 20194
rect 435548 20130 435600 20136
rect 435364 17468 435416 17474
rect 435364 17410 435416 17416
rect 435560 13870 435588 20130
rect 437480 19440 437532 19446
rect 437480 19382 437532 19388
rect 436008 17604 436060 17610
rect 436008 17546 436060 17552
rect 435824 14816 435876 14822
rect 435824 14758 435876 14764
rect 435548 13864 435600 13870
rect 435548 13806 435600 13812
rect 432052 13456 432104 13462
rect 432052 13398 432104 13404
rect 431408 11756 431460 11762
rect 431408 11698 431460 11704
rect 430580 9036 430632 9042
rect 430580 8978 430632 8984
rect 431316 9036 431368 9042
rect 431316 8978 431368 8984
rect 428462 7984 428518 7993
rect 428462 7919 428518 7928
rect 427728 6656 427780 6662
rect 427728 6598 427780 6604
rect 426900 6384 426952 6390
rect 426900 6326 426952 6332
rect 427176 6384 427228 6390
rect 427176 6326 427228 6332
rect 426162 3632 426218 3641
rect 426162 3567 426218 3576
rect 426176 480 426204 3567
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426912 354 426940 6326
rect 427728 6316 427780 6322
rect 427728 6258 427780 6264
rect 427740 2854 427768 6258
rect 427728 2848 427780 2854
rect 427728 2790 427780 2796
rect 428476 480 428504 7919
rect 430592 3738 430620 8978
rect 431420 6798 431448 11698
rect 431408 6792 431460 6798
rect 431408 6734 431460 6740
rect 430856 6588 430908 6594
rect 430856 6530 430908 6536
rect 430580 3732 430632 3738
rect 430580 3674 430632 3680
rect 429660 2848 429712 2854
rect 429660 2790 429712 2796
rect 429672 480 429700 2790
rect 430868 480 430896 6530
rect 432064 480 432092 13398
rect 433984 12300 434036 12306
rect 433984 12242 434036 12248
rect 433996 6594 434024 12242
rect 434904 12028 434956 12034
rect 434904 11970 434956 11976
rect 434916 9654 434944 11970
rect 435836 11898 435864 14758
rect 436020 12374 436048 17546
rect 437492 16862 437520 19382
rect 438124 17332 438176 17338
rect 438124 17274 438176 17280
rect 437480 16856 437532 16862
rect 437480 16798 437532 16804
rect 436744 16176 436796 16182
rect 436744 16118 436796 16124
rect 435916 12368 435968 12374
rect 435916 12310 435968 12316
rect 436008 12368 436060 12374
rect 436008 12310 436060 12316
rect 435824 11892 435876 11898
rect 435824 11834 435876 11840
rect 434904 9648 434956 9654
rect 434904 9590 434956 9596
rect 435928 9246 435956 12310
rect 435456 9240 435508 9246
rect 435456 9182 435508 9188
rect 435916 9240 435968 9246
rect 435916 9182 435968 9188
rect 434628 6792 434680 6798
rect 434628 6734 434680 6740
rect 433984 6588 434036 6594
rect 433984 6530 434036 6536
rect 434444 3732 434496 3738
rect 434444 3674 434496 3680
rect 433248 3596 433300 3602
rect 433248 3538 433300 3544
rect 433260 480 433288 3538
rect 434456 480 434484 3674
rect 434640 3194 434668 6734
rect 435468 6322 435496 9182
rect 436008 9172 436060 9178
rect 436008 9114 436060 9120
rect 435456 6316 435508 6322
rect 435456 6258 435508 6264
rect 435546 6216 435602 6225
rect 435546 6151 435602 6160
rect 434628 3188 434680 3194
rect 434628 3130 434680 3136
rect 435560 480 435588 6151
rect 436020 3602 436048 9114
rect 436008 3596 436060 3602
rect 436008 3538 436060 3544
rect 436756 480 436784 16118
rect 438136 9382 438164 17274
rect 438872 17066 438900 22238
rect 439516 20194 439544 154119
rect 439504 20188 439556 20194
rect 439504 20130 439556 20136
rect 439228 18896 439280 18902
rect 439228 18838 439280 18844
rect 438860 17060 438912 17066
rect 438860 17002 438912 17008
rect 438860 16108 438912 16114
rect 438860 16050 438912 16056
rect 438872 11762 438900 16050
rect 439240 14822 439268 18838
rect 442276 17950 442304 155071
rect 442264 17944 442316 17950
rect 442264 17886 442316 17892
rect 439412 17536 439464 17542
rect 439412 17478 439464 17484
rect 439424 14958 439452 17478
rect 441988 17060 442040 17066
rect 441988 17002 442040 17008
rect 441620 16856 441672 16862
rect 441620 16798 441672 16804
rect 439412 14952 439464 14958
rect 439412 14894 439464 14900
rect 439228 14816 439280 14822
rect 439228 14758 439280 14764
rect 440884 13864 440936 13870
rect 440884 13806 440936 13812
rect 440240 11960 440292 11966
rect 440240 11902 440292 11908
rect 438860 11756 438912 11762
rect 438860 11698 438912 11704
rect 438768 9648 438820 9654
rect 438768 9590 438820 9596
rect 438124 9376 438176 9382
rect 438124 9318 438176 9324
rect 438780 3670 438808 9590
rect 440252 9314 440280 11902
rect 440240 9308 440292 9314
rect 440240 9250 440292 9256
rect 439134 5128 439190 5137
rect 439134 5063 439190 5072
rect 438768 3664 438820 3670
rect 438768 3606 438820 3612
rect 437940 3188 437992 3194
rect 437940 3130 437992 3136
rect 437952 480 437980 3130
rect 439148 480 439176 5063
rect 440896 3602 440924 13806
rect 441632 12442 441660 16798
rect 442000 14278 442028 17002
rect 442908 14952 442960 14958
rect 442908 14894 442960 14900
rect 441988 14272 442040 14278
rect 441988 14214 442040 14220
rect 441620 12436 441672 12442
rect 441620 12378 441672 12384
rect 442920 12306 442948 14894
rect 445036 14414 445064 160142
rect 445760 25084 445812 25090
rect 445760 25026 445812 25032
rect 445484 17944 445536 17950
rect 445484 17886 445536 17892
rect 445116 14816 445168 14822
rect 445116 14758 445168 14764
rect 445024 14408 445076 14414
rect 445024 14350 445076 14356
rect 444656 12436 444708 12442
rect 444656 12378 444708 12384
rect 442908 12300 442960 12306
rect 442908 12242 442960 12248
rect 443368 12232 443420 12238
rect 443368 12174 443420 12180
rect 442630 10296 442686 10305
rect 442630 10231 442686 10240
rect 441528 6656 441580 6662
rect 441528 6598 441580 6604
rect 440332 3596 440384 3602
rect 440332 3538 440384 3544
rect 440884 3596 440936 3602
rect 440884 3538 440936 3544
rect 440344 480 440372 3538
rect 441540 480 441568 6598
rect 442644 480 442672 10231
rect 427238 354 427350 480
rect 426912 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 12174
rect 444668 8430 444696 12378
rect 445024 9036 445076 9042
rect 445024 8978 445076 8984
rect 444656 8424 444708 8430
rect 444656 8366 444708 8372
rect 445036 480 445064 8978
rect 445128 3126 445156 14758
rect 445496 11694 445524 17886
rect 445668 11756 445720 11762
rect 445668 11698 445720 11704
rect 445484 11688 445536 11694
rect 445484 11630 445536 11636
rect 445680 9042 445708 11698
rect 445668 9036 445720 9042
rect 445668 8978 445720 8984
rect 445116 3120 445168 3126
rect 445116 3062 445168 3068
rect 445668 2848 445720 2854
rect 445668 2790 445720 2796
rect 445680 2718 445708 2790
rect 445668 2712 445720 2718
rect 445668 2654 445720 2660
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 25026
rect 448704 17468 448756 17474
rect 448704 17410 448756 17416
rect 448716 14822 448744 17410
rect 449176 14958 449204 161502
rect 463700 160132 463752 160138
rect 463700 160074 463752 160080
rect 454684 157412 454736 157418
rect 454684 157354 454736 157360
rect 453304 152040 453356 152046
rect 453304 151982 453356 151988
rect 453316 23186 453344 151982
rect 453304 23180 453356 23186
rect 453304 23122 453356 23128
rect 453304 20188 453356 20194
rect 453304 20130 453356 20136
rect 449164 14952 449216 14958
rect 449164 14894 449216 14900
rect 448704 14816 448756 14822
rect 448704 14758 448756 14764
rect 450912 14748 450964 14754
rect 450912 14690 450964 14696
rect 448520 14408 448572 14414
rect 448520 14350 448572 14356
rect 448532 12102 448560 14350
rect 448612 14272 448664 14278
rect 448612 14214 448664 14220
rect 448520 12096 448572 12102
rect 448520 12038 448572 12044
rect 448624 11966 448652 14214
rect 449808 12368 449860 12374
rect 449808 12310 449860 12316
rect 448796 12300 448848 12306
rect 448796 12242 448848 12248
rect 448808 12034 448836 12242
rect 448704 12028 448756 12034
rect 448704 11970 448756 11976
rect 448796 12028 448848 12034
rect 448796 11970 448848 11976
rect 448612 11960 448664 11966
rect 448612 11902 448664 11908
rect 448716 9178 448744 11970
rect 449164 10464 449216 10470
rect 449164 10406 449216 10412
rect 448704 9172 448756 9178
rect 448704 9114 448756 9120
rect 449176 6730 449204 10406
rect 449440 9376 449492 9382
rect 449440 9318 449492 9324
rect 449164 6724 449216 6730
rect 449164 6666 449216 6672
rect 448520 6588 448572 6594
rect 448520 6530 448572 6536
rect 448532 3874 448560 6530
rect 449452 6526 449480 9318
rect 449820 9194 449848 12310
rect 449820 9166 449940 9194
rect 449912 9110 449940 9166
rect 449808 9104 449860 9110
rect 449808 9046 449860 9052
rect 449900 9104 449952 9110
rect 449900 9046 449952 9052
rect 448612 6520 448664 6526
rect 448612 6462 448664 6468
rect 449440 6520 449492 6526
rect 449440 6462 449492 6468
rect 448520 3868 448572 3874
rect 448520 3810 448572 3816
rect 448624 3738 448652 6462
rect 448612 3732 448664 3738
rect 448612 3674 448664 3680
rect 448612 3120 448664 3126
rect 448612 3062 448664 3068
rect 447416 2848 447468 2854
rect 447416 2790 447468 2796
rect 447428 480 447456 2790
rect 448624 480 448652 3062
rect 449820 480 449848 9046
rect 450924 480 450952 14690
rect 453316 11694 453344 20130
rect 453304 11688 453356 11694
rect 453210 11656 453266 11665
rect 453304 11630 453356 11636
rect 453210 11591 453266 11600
rect 452752 9308 452804 9314
rect 452752 9250 452804 9256
rect 452660 8424 452712 8430
rect 452660 8366 452712 8372
rect 452672 3806 452700 8366
rect 452660 3800 452712 3806
rect 452660 3742 452712 3748
rect 452764 3602 452792 9250
rect 453224 6914 453252 11591
rect 453224 6886 453344 6914
rect 452108 3596 452160 3602
rect 452108 3538 452160 3544
rect 452752 3596 452804 3602
rect 452752 3538 452804 3544
rect 452120 480 452148 3538
rect 453316 480 453344 6886
rect 454696 5574 454724 157354
rect 462964 153400 463016 153406
rect 462964 153342 463016 153348
rect 458824 151972 458876 151978
rect 458824 151914 458876 151920
rect 458180 23180 458232 23186
rect 458180 23122 458232 23128
rect 458192 20194 458220 23122
rect 458180 20188 458232 20194
rect 458180 20130 458232 20136
rect 454776 17400 454828 17406
rect 454776 17342 454828 17348
rect 454788 5642 454816 17342
rect 456064 14952 456116 14958
rect 456064 14894 456116 14900
rect 456076 9314 456104 14894
rect 457444 11688 457496 11694
rect 457444 11630 457496 11636
rect 456064 9308 456116 9314
rect 456064 9250 456116 9256
rect 455696 6724 455748 6730
rect 455696 6666 455748 6672
rect 454776 5636 454828 5642
rect 454776 5578 454828 5584
rect 454684 5568 454736 5574
rect 454684 5510 454736 5516
rect 454498 3496 454554 3505
rect 454498 3431 454554 3440
rect 454512 480 454540 3431
rect 455708 480 455736 6666
rect 457456 3602 457484 11630
rect 458836 9246 458864 151914
rect 460204 151904 460256 151910
rect 460204 151846 460256 151852
rect 459192 12028 459244 12034
rect 459192 11970 459244 11976
rect 458088 9240 458140 9246
rect 458088 9182 458140 9188
rect 458824 9240 458876 9246
rect 458824 9182 458876 9188
rect 458100 6594 458128 9182
rect 458088 6588 458140 6594
rect 458088 6530 458140 6536
rect 458088 6452 458140 6458
rect 458088 6394 458140 6400
rect 456892 3596 456944 3602
rect 456892 3538 456944 3544
rect 457444 3596 457496 3602
rect 457444 3538 457496 3544
rect 456904 480 456932 3538
rect 458100 480 458128 6394
rect 459204 480 459232 11970
rect 460216 6458 460244 151846
rect 462976 23458 463004 153342
rect 462964 23452 463016 23458
rect 462964 23394 463016 23400
rect 460296 19508 460348 19514
rect 460296 19450 460348 19456
rect 460308 14754 460336 19450
rect 463712 16574 463740 160074
rect 494072 156670 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 162081 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 527178 162072 527234 162081
rect 527178 162007 527234 162016
rect 557540 161492 557592 161498
rect 557540 161434 557592 161440
rect 494060 156664 494112 156670
rect 494060 156606 494112 156612
rect 529940 155644 529992 155650
rect 529940 155586 529992 155592
rect 507858 155000 507914 155009
rect 507858 154935 507914 154944
rect 485044 153876 485096 153882
rect 485044 153818 485096 153824
rect 485056 152522 485084 153818
rect 489920 153332 489972 153338
rect 489920 153274 489972 153280
rect 485044 152516 485096 152522
rect 485044 152458 485096 152464
rect 467104 152312 467156 152318
rect 467104 152254 467156 152260
rect 466736 23452 466788 23458
rect 466736 23394 466788 23400
rect 466748 20670 466776 23394
rect 466736 20664 466788 20670
rect 466736 20606 466788 20612
rect 463712 16546 464016 16574
rect 460296 14748 460348 14754
rect 460296 14690 460348 14696
rect 463148 12164 463200 12170
rect 463148 12106 463200 12112
rect 460296 12096 460348 12102
rect 460296 12038 460348 12044
rect 460204 6452 460256 6458
rect 460204 6394 460256 6400
rect 459560 5636 459612 5642
rect 459560 5578 459612 5584
rect 459572 3942 459600 5578
rect 460308 4010 460336 12038
rect 463160 9518 463188 12106
rect 463148 9512 463200 9518
rect 463148 9454 463200 9460
rect 462318 9072 462374 9081
rect 462318 9007 462374 9016
rect 462332 6730 462360 9007
rect 462320 6724 462372 6730
rect 462320 6666 462372 6672
rect 462504 6384 462556 6390
rect 462504 6326 462556 6332
rect 460296 4004 460348 4010
rect 460296 3946 460348 3952
rect 459560 3936 459612 3942
rect 459560 3878 459612 3884
rect 462516 3670 462544 6326
rect 462780 5568 462832 5574
rect 462780 5510 462832 5516
rect 460388 3664 460440 3670
rect 460388 3606 460440 3612
rect 462504 3664 462556 3670
rect 462504 3606 462556 3612
rect 460400 480 460428 3606
rect 461582 3360 461638 3369
rect 461582 3295 461638 3304
rect 461596 480 461624 3295
rect 462792 480 462820 5510
rect 463988 480 464016 16546
rect 467116 6662 467144 152254
rect 476764 151496 476816 151502
rect 476764 151438 476816 151444
rect 471428 22772 471480 22778
rect 471428 22714 471480 22720
rect 471336 20664 471388 20670
rect 471336 20606 471388 20612
rect 467196 20188 467248 20194
rect 467196 20130 467248 20136
rect 467104 6656 467156 6662
rect 467104 6598 467156 6604
rect 467208 6526 467236 20130
rect 470600 18828 470652 18834
rect 470600 18770 470652 18776
rect 470612 12034 470640 18770
rect 471348 17950 471376 20606
rect 471336 17944 471388 17950
rect 471336 17886 471388 17892
rect 471440 17882 471468 22714
rect 474004 17944 474056 17950
rect 474004 17886 474056 17892
rect 471428 17876 471480 17882
rect 471428 17818 471480 17824
rect 471980 17264 472032 17270
rect 471980 17206 472032 17212
rect 471992 16574 472020 17206
rect 471992 16546 472296 16574
rect 471244 14748 471296 14754
rect 471244 14690 471296 14696
rect 470600 12028 470652 12034
rect 470600 11970 470652 11976
rect 467656 9512 467708 9518
rect 467656 9454 467708 9460
rect 467564 6588 467616 6594
rect 467564 6530 467616 6536
rect 465172 6520 465224 6526
rect 465172 6462 465224 6468
rect 467196 6520 467248 6526
rect 467196 6462 467248 6468
rect 465184 480 465212 6462
rect 466460 6248 466512 6254
rect 466460 6190 466512 6196
rect 466472 3806 466500 6190
rect 467576 3942 467604 6530
rect 467668 6390 467696 9454
rect 470692 9240 470744 9246
rect 470692 9182 470744 9188
rect 467656 6384 467708 6390
rect 467656 6326 467708 6332
rect 470704 6254 470732 9182
rect 471060 6724 471112 6730
rect 471060 6666 471112 6672
rect 470692 6248 470744 6254
rect 470692 6190 470744 6196
rect 469864 4004 469916 4010
rect 469864 3946 469916 3952
rect 467472 3936 467524 3942
rect 467472 3878 467524 3884
rect 467564 3936 467616 3942
rect 467564 3878 467616 3884
rect 466276 3800 466328 3806
rect 466276 3742 466328 3748
rect 466460 3800 466512 3806
rect 466460 3742 466512 3748
rect 466288 480 466316 3742
rect 467484 480 467512 3878
rect 468668 3528 468720 3534
rect 468668 3470 468720 3476
rect 468680 480 468708 3470
rect 469876 480 469904 3946
rect 471072 480 471100 6666
rect 471256 5574 471284 14690
rect 471980 9308 472032 9314
rect 471980 9250 472032 9256
rect 471992 6730 472020 9250
rect 471980 6724 472032 6730
rect 471980 6666 472032 6672
rect 471888 6316 471940 6322
rect 471888 6258 471940 6264
rect 471244 5568 471296 5574
rect 471244 5510 471296 5516
rect 471900 3262 471928 6258
rect 471888 3256 471940 3262
rect 471888 3198 471940 3204
rect 472268 480 472296 16546
rect 474016 9314 474044 17886
rect 475384 17876 475436 17882
rect 475384 17818 475436 17824
rect 474004 9308 474056 9314
rect 474004 9250 474056 9256
rect 475396 6458 475424 17818
rect 476776 17134 476804 151438
rect 485044 25560 485096 25566
rect 485044 25502 485096 25508
rect 480904 22840 480956 22846
rect 480904 22782 480956 22788
rect 477408 17672 477460 17678
rect 477408 17614 477460 17620
rect 476764 17128 476816 17134
rect 476764 17070 476816 17076
rect 476764 16040 476816 16046
rect 476764 15982 476816 15988
rect 476028 9172 476080 9178
rect 476028 9114 476080 9120
rect 476040 6798 476068 9114
rect 476028 6792 476080 6798
rect 476028 6734 476080 6740
rect 476776 6594 476804 15982
rect 477420 14890 477448 17614
rect 480260 17128 480312 17134
rect 480260 17070 480312 17076
rect 478144 15972 478196 15978
rect 478144 15914 478196 15920
rect 477408 14884 477460 14890
rect 477408 14826 477460 14832
rect 476764 6588 476816 6594
rect 476764 6530 476816 6536
rect 473820 6452 473872 6458
rect 473820 6394 473872 6400
rect 475384 6452 475436 6458
rect 475384 6394 475436 6400
rect 473832 3534 473860 6394
rect 476948 5568 477000 5574
rect 476948 5510 477000 5516
rect 474556 3868 474608 3874
rect 474556 3810 474608 3816
rect 473820 3528 473872 3534
rect 473820 3470 473872 3476
rect 473452 3256 473504 3262
rect 473452 3198 473504 3204
rect 473464 480 473492 3198
rect 474568 480 474596 3810
rect 475752 3460 475804 3466
rect 475752 3402 475804 3408
rect 475764 480 475792 3402
rect 476960 480 476988 5510
rect 478156 480 478184 15914
rect 480272 14754 480300 17070
rect 480260 14748 480312 14754
rect 480260 14690 480312 14696
rect 480916 11694 480944 22782
rect 482374 13016 482430 13025
rect 482374 12951 482430 12960
rect 480904 11688 480956 11694
rect 480904 11630 480956 11636
rect 478880 9036 478932 9042
rect 478880 8978 478932 8984
rect 478892 6322 478920 8978
rect 481732 6724 481784 6730
rect 481732 6666 481784 6672
rect 480536 6656 480588 6662
rect 480536 6598 480588 6604
rect 478880 6316 478932 6322
rect 478880 6258 478932 6264
rect 479340 3936 479392 3942
rect 479340 3878 479392 3884
rect 479352 480 479380 3878
rect 480548 480 480576 6598
rect 481548 6248 481600 6254
rect 481548 6190 481600 6196
rect 481560 3194 481588 6190
rect 481548 3188 481600 3194
rect 481548 3130 481600 3136
rect 481744 480 481772 6666
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 12951
rect 485056 12102 485084 25502
rect 488540 25016 488592 25022
rect 488540 24958 488592 24964
rect 488552 16574 488580 24958
rect 489932 16574 489960 153274
rect 503720 151224 503772 151230
rect 503720 151166 503772 151172
rect 491944 151156 491996 151162
rect 491944 151098 491996 151104
rect 488552 16546 488856 16574
rect 489932 16546 490696 16574
rect 485136 15904 485188 15910
rect 485136 15846 485188 15852
rect 485044 12096 485096 12102
rect 485044 12038 485096 12044
rect 484860 6792 484912 6798
rect 484860 6734 484912 6740
rect 484400 6520 484452 6526
rect 484400 6462 484452 6468
rect 484412 3330 484440 6462
rect 484400 3324 484452 3330
rect 484400 3266 484452 3272
rect 484032 3188 484084 3194
rect 484032 3130 484084 3136
rect 484044 480 484072 3130
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484872 354 484900 6734
rect 485148 6526 485176 15846
rect 488632 14884 488684 14890
rect 488632 14826 488684 14832
rect 488644 11898 488672 14826
rect 488540 11892 488592 11898
rect 488540 11834 488592 11840
rect 488632 11892 488684 11898
rect 488632 11834 488684 11840
rect 485228 11688 485280 11694
rect 485228 11630 485280 11636
rect 485136 6520 485188 6526
rect 485136 6462 485188 6468
rect 485240 6254 485268 11630
rect 488552 9178 488580 11834
rect 488540 9172 488592 9178
rect 488540 9114 488592 9120
rect 486422 7848 486478 7857
rect 486422 7783 486478 7792
rect 485228 6248 485280 6254
rect 485228 6190 485280 6196
rect 486436 480 486464 7783
rect 487620 3324 487672 3330
rect 487620 3266 487672 3272
rect 487632 480 487660 3266
rect 488828 480 488856 16546
rect 489920 4888 489972 4894
rect 489920 4830 489972 4836
rect 489932 480 489960 4830
rect 485198 354 485310 480
rect 484872 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 491208 11960 491260 11966
rect 491208 11902 491260 11908
rect 491220 9382 491248 11902
rect 491208 9376 491260 9382
rect 491208 9318 491260 9324
rect 491300 9308 491352 9314
rect 491300 9250 491352 9256
rect 491312 5574 491340 9250
rect 491956 9246 491984 151098
rect 494704 24948 494756 24954
rect 494704 24890 494756 24896
rect 494716 16574 494744 24890
rect 495440 20120 495492 20126
rect 495440 20062 495492 20068
rect 494716 16546 494836 16574
rect 493324 14680 493376 14686
rect 493324 14622 493376 14628
rect 491944 9240 491996 9246
rect 491944 9182 491996 9188
rect 492312 6588 492364 6594
rect 492312 6530 492364 6536
rect 492036 6384 492088 6390
rect 492036 6326 492088 6332
rect 491300 5568 491352 5574
rect 491300 5510 491352 5516
rect 492048 3466 492076 6326
rect 492036 3460 492088 3466
rect 492036 3402 492088 3408
rect 492324 480 492352 6530
rect 493336 6390 493364 14622
rect 493968 11892 494020 11898
rect 493968 11834 494020 11840
rect 493980 9042 494008 11834
rect 493968 9036 494020 9042
rect 493968 8978 494020 8984
rect 493508 6520 493560 6526
rect 493508 6462 493560 6468
rect 493324 6384 493376 6390
rect 493324 6326 493376 6332
rect 493520 480 493548 6462
rect 494704 5568 494756 5574
rect 494704 5510 494756 5516
rect 494716 480 494744 5510
rect 494808 3874 494836 16546
rect 494796 3868 494848 3874
rect 494796 3810 494848 3816
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 354 495480 20062
rect 499580 20052 499632 20058
rect 499580 19994 499632 20000
rect 499592 16574 499620 19994
rect 502984 18624 503036 18630
rect 502984 18566 503036 18572
rect 499592 16546 500632 16574
rect 498936 14544 498988 14550
rect 498936 14486 498988 14492
rect 498292 12096 498344 12102
rect 498292 12038 498344 12044
rect 498304 9110 498332 12038
rect 498200 9104 498252 9110
rect 498200 9046 498252 9052
rect 498292 9104 498344 9110
rect 498292 9046 498344 9052
rect 497096 3800 497148 3806
rect 497096 3742 497148 3748
rect 497108 480 497136 3742
rect 498212 480 498240 9046
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 14486
rect 500604 480 500632 16546
rect 502996 9654 503024 18566
rect 502984 9648 503036 9654
rect 502984 9590 503036 9596
rect 503628 8968 503680 8974
rect 503628 8910 503680 8916
rect 502984 6452 503036 6458
rect 502984 6394 503036 6400
rect 501788 3528 501840 3534
rect 501788 3470 501840 3476
rect 501800 480 501828 3470
rect 502996 480 503024 6394
rect 503640 3534 503668 8910
rect 503628 3528 503680 3534
rect 503628 3470 503680 3476
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 151166
rect 507124 20868 507176 20874
rect 507124 20810 507176 20816
rect 506480 9648 506532 9654
rect 506480 9590 506532 9596
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 505388 480 505416 3470
rect 506492 480 506520 9590
rect 507136 9314 507164 20810
rect 507872 16574 507900 154935
rect 512642 154864 512698 154873
rect 512642 154799 512698 154808
rect 509884 26376 509936 26382
rect 509884 26318 509936 26324
rect 507872 16546 508912 16574
rect 507216 14748 507268 14754
rect 507216 14690 507268 14696
rect 507124 9308 507176 9314
rect 507124 9250 507176 9256
rect 507228 6866 507256 14690
rect 507216 6860 507268 6866
rect 507216 6802 507268 6808
rect 507676 3868 507728 3874
rect 507676 3810 507728 3816
rect 507688 480 507716 3810
rect 508884 480 508912 16546
rect 509608 6860 509660 6866
rect 509608 6802 509660 6808
rect 509620 3534 509648 6802
rect 509896 6594 509924 26318
rect 510620 26308 510672 26314
rect 510620 26250 510672 26256
rect 510632 16574 510660 26250
rect 510632 16546 511304 16574
rect 510252 12028 510304 12034
rect 510252 11970 510304 11976
rect 510264 9450 510292 11970
rect 510252 9444 510304 9450
rect 510252 9386 510304 9392
rect 510068 9376 510120 9382
rect 510068 9318 510120 9324
rect 509884 6588 509936 6594
rect 509884 6530 509936 6536
rect 509608 3528 509660 3534
rect 509608 3470 509660 3476
rect 510080 480 510108 9318
rect 511276 480 511304 16546
rect 512000 11756 512052 11762
rect 512000 11698 512052 11704
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 11698
rect 512656 3194 512684 154799
rect 525800 153264 525852 153270
rect 525800 153206 525852 153212
rect 516784 152516 516836 152522
rect 516784 152458 516836 152464
rect 513380 19372 513432 19378
rect 513380 19314 513432 19320
rect 513288 14816 513340 14822
rect 513288 14758 513340 14764
rect 513300 11762 513328 14758
rect 513288 11756 513340 11762
rect 513288 11698 513340 11704
rect 512644 3188 512696 3194
rect 512644 3130 512696 3136
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 19314
rect 516140 13116 516192 13122
rect 516140 13058 516192 13064
rect 516152 8974 516180 13058
rect 516140 8968 516192 8974
rect 516140 8910 516192 8916
rect 516796 4146 516824 152458
rect 525812 16574 525840 153206
rect 527178 19408 527234 19417
rect 527178 19343 527234 19352
rect 527192 16574 527220 19343
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 521660 14612 521712 14618
rect 521660 14554 521712 14560
rect 520280 13252 520332 13258
rect 520280 13194 520332 13200
rect 517152 9444 517204 9450
rect 517152 9386 517204 9392
rect 516784 4140 516836 4146
rect 516784 4082 516836 4088
rect 514760 3732 514812 3738
rect 514760 3674 514812 3680
rect 514772 480 514800 3674
rect 515956 3188 516008 3194
rect 515956 3130 516008 3136
rect 515968 480 515996 3130
rect 517164 480 517192 9386
rect 518346 7712 518402 7721
rect 518346 7647 518402 7656
rect 518360 480 518388 7647
rect 519544 4140 519596 4146
rect 519544 4082 519596 4088
rect 519556 480 519584 4082
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 13194
rect 520924 11824 520976 11830
rect 520924 11766 520976 11772
rect 520936 6458 520964 11766
rect 520924 6452 520976 6458
rect 520924 6394 520976 6400
rect 521568 4820 521620 4826
rect 521568 4762 521620 4768
rect 521580 2854 521608 4762
rect 521568 2848 521620 2854
rect 521568 2790 521620 2796
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 14554
rect 525800 6384 525852 6390
rect 525800 6326 525852 6332
rect 525430 4992 525486 5001
rect 525430 4927 525486 4936
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523052 480 523080 3470
rect 524236 2848 524288 2854
rect 524236 2790 524288 2796
rect 524248 480 524276 2790
rect 525444 480 525472 4927
rect 525812 3534 525840 6326
rect 525800 3528 525852 3534
rect 525800 3470 525852 3476
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 526260 9172 526312 9178
rect 526260 9114 526312 9120
rect 526272 6390 526300 9114
rect 526260 6384 526312 6390
rect 526260 6326 526312 6332
rect 527836 480 527864 16546
rect 528560 9240 528612 9246
rect 528560 9182 528612 9188
rect 528572 6526 528600 9182
rect 529020 6588 529072 6594
rect 529020 6530 529072 6536
rect 528560 6520 528612 6526
rect 528560 6462 528612 6468
rect 529032 480 529060 6530
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 529952 354 529980 155586
rect 539598 154728 539654 154737
rect 539598 154663 539654 154672
rect 534724 20800 534776 20806
rect 534724 20742 534776 20748
rect 532056 15224 532108 15230
rect 532056 15166 532108 15172
rect 531228 11756 531280 11762
rect 531228 11698 531280 11704
rect 531240 9178 531268 11698
rect 531228 9172 531280 9178
rect 531228 9114 531280 9120
rect 531320 9104 531372 9110
rect 531320 9046 531372 9052
rect 531332 480 531360 9046
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 15166
rect 534736 9110 534764 20742
rect 539612 16574 539640 154663
rect 543738 152144 543794 152153
rect 543738 152079 543794 152088
rect 542360 19984 542412 19990
rect 542360 19926 542412 19932
rect 542372 16574 542400 19926
rect 543752 16574 543780 152079
rect 556160 24880 556212 24886
rect 556160 24822 556212 24828
rect 549260 24132 549312 24138
rect 549260 24074 549312 24080
rect 545118 18592 545174 18601
rect 545118 18527 545174 18536
rect 545132 16574 545160 18527
rect 549272 16574 549300 24074
rect 553400 23724 553452 23730
rect 553400 23666 553452 23672
rect 552020 20732 552072 20738
rect 552020 20674 552072 20680
rect 552032 16574 552060 20674
rect 553412 16574 553440 23666
rect 556172 16574 556200 24822
rect 557552 16574 557580 161434
rect 558932 156641 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 579908 218074 579936 218991
rect 579896 218068 579948 218074
rect 579896 218010 579948 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580276 158001 580304 670647
rect 580262 157992 580318 158001
rect 580262 157927 580318 157936
rect 558918 156632 558974 156641
rect 558918 156567 558974 156576
rect 576122 154592 576178 154601
rect 576122 154527 576178 154536
rect 561680 151088 561732 151094
rect 561680 151030 561732 151036
rect 560300 18692 560352 18698
rect 560300 18634 560352 18640
rect 560312 16574 560340 18634
rect 561692 16574 561720 151030
rect 576136 60722 576164 154527
rect 578884 153468 578936 153474
rect 578884 153410 578936 153416
rect 576124 60716 576176 60722
rect 576124 60658 576176 60664
rect 563060 23656 563112 23662
rect 563060 23598 563112 23604
rect 539612 16546 540376 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 534816 10328 534868 10334
rect 534816 10270 534868 10276
rect 534724 9104 534776 9110
rect 534724 9046 534776 9052
rect 534828 5574 534856 10270
rect 534908 9308 534960 9314
rect 534908 9250 534960 9256
rect 534816 5568 534868 5574
rect 534816 5510 534868 5516
rect 533712 3664 533764 3670
rect 533712 3606 533764 3612
rect 533724 480 533752 3606
rect 534920 480 534948 9250
rect 538402 8936 538458 8945
rect 538402 8871 538458 8880
rect 536104 6180 536156 6186
rect 536104 6122 536156 6128
rect 536116 480 536144 6122
rect 537208 3596 537260 3602
rect 537208 3538 537260 3544
rect 537220 480 537248 3538
rect 538416 480 538444 8871
rect 539600 5568 539652 5574
rect 539600 5510 539652 5516
rect 539612 480 539640 5510
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 9172 542044 9178
rect 541992 9114 542044 9120
rect 542004 480 542032 9114
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543740 6316 543792 6322
rect 543740 6258 543792 6264
rect 543752 3602 543780 6258
rect 543740 3596 543792 3602
rect 543740 3538 543792 3544
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 548616 10396 548668 10402
rect 548616 10338 548668 10344
rect 547880 6520 547932 6526
rect 547880 6462 547932 6468
rect 546684 6452 546736 6458
rect 546684 6394 546736 6400
rect 546696 480 546724 6394
rect 547892 480 547920 6462
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 10338
rect 550284 480 550312 16546
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 551480 480 551508 3538
rect 552572 2848 552624 2854
rect 552572 2790 552624 2796
rect 552584 2689 552612 2790
rect 552570 2680 552626 2689
rect 552570 2615 552626 2624
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554964 3528 555016 3534
rect 554964 3470 555016 3476
rect 554976 480 555004 3470
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 82 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 559748 2848 559800 2854
rect 559748 2790 559800 2796
rect 559760 480 559788 2790
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 556342 96 556398 105
rect 556130 54 556342 82
rect 556130 -960 556242 54
rect 556342 31 556398 40
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 562322 7576 562378 7585
rect 562322 7511 562378 7520
rect 562336 3534 562364 7511
rect 562324 3528 562376 3534
rect 562324 3470 562376 3476
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 23598
rect 571340 23588 571392 23594
rect 571340 23530 571392 23536
rect 567200 22228 567252 22234
rect 567200 22170 567252 22176
rect 567212 16574 567240 22170
rect 567212 16546 567608 16574
rect 565820 9036 565872 9042
rect 565820 8978 565872 8984
rect 565636 6384 565688 6390
rect 565636 6326 565688 6332
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564452 480 564480 3470
rect 565648 480 565676 6326
rect 565832 3330 565860 8978
rect 566832 6248 566884 6254
rect 566832 6190 566884 6196
rect 565820 3324 565872 3330
rect 565820 3266 565872 3272
rect 566844 480 566872 6190
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 570328 14476 570380 14482
rect 570328 14418 570380 14424
rect 569132 3324 569184 3330
rect 569132 3266 569184 3272
rect 569144 480 569172 3266
rect 570340 480 570368 14418
rect 571248 9104 571300 9110
rect 571248 9046 571300 9052
rect 571260 3534 571288 9046
rect 571248 3528 571300 3534
rect 571248 3470 571300 3476
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 23530
rect 575480 23520 575532 23526
rect 575480 23462 575532 23468
rect 574100 22160 574152 22166
rect 574100 22102 574152 22108
rect 574112 16574 574140 22102
rect 575492 16574 575520 23462
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 572720 2848 572772 2854
rect 572720 2790 572772 2796
rect 572732 480 572760 2790
rect 573928 480 573956 3470
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 577424 480 577452 8910
rect 578896 6633 578924 153410
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580276 19825 580304 152623
rect 582378 24984 582434 24993
rect 582378 24919 582434 24928
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 581090 17232 581146 17241
rect 581090 17167 581146 17176
rect 581104 16574 581132 17167
rect 582392 16574 582420 24919
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 578882 6624 578938 6633
rect 578882 6559 578938 6568
rect 578606 4856 578662 4865
rect 578606 4791 578662 4800
rect 578620 480 578648 4791
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3146 214920 3202 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3422 162868 3424 162888
rect 3424 162868 3476 162888
rect 3476 162868 3478 162888
rect 3422 162832 3478 162868
rect 3422 149776 3478 149832
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3146 97552 3202 97608
rect 2962 84632 3018 84688
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 3330 58520 3386 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 3146 19352 3202 19408
rect 3514 6432 3570 6488
rect 9126 160112 9182 160168
rect 9494 15136 9550 15192
rect 10506 151816 10562 151872
rect 13174 16632 13230 16688
rect 12346 12960 12402 13016
rect 10966 9560 11022 9616
rect 13634 153720 13690 153776
rect 13542 153176 13598 153232
rect 14462 156032 14518 156088
rect 14554 153312 14610 153368
rect 14830 154672 14886 154728
rect 14738 154128 14794 154184
rect 14830 16496 14886 16552
rect 14738 15816 14794 15872
rect 15014 14456 15070 14512
rect 16026 19896 16082 19952
rect 18050 159296 18106 159352
rect 18234 157392 18290 157448
rect 17682 18672 17738 18728
rect 17406 18536 17462 18592
rect 17682 17720 17738 17776
rect 18878 17856 18934 17912
rect 19154 154944 19210 155000
rect 18970 17176 19026 17232
rect 18694 16632 18750 16688
rect 19706 155080 19762 155136
rect 19798 154808 19854 154864
rect 19154 12280 19210 12336
rect 19706 19216 19762 19272
rect 20166 16224 20222 16280
rect 20626 158752 20682 158808
rect 22098 155352 22154 155408
rect 22098 153720 22154 153776
rect 26146 153720 26202 153776
rect 22190 153584 22246 153640
rect 24306 153448 24362 153504
rect 25410 152632 25466 152688
rect 28722 154536 28778 154592
rect 35622 155352 35678 155408
rect 31666 155216 31722 155272
rect 28906 154400 28962 154456
rect 29826 153856 29882 153912
rect 30838 153584 30894 153640
rect 33046 152496 33102 152552
rect 34978 153992 35034 154048
rect 35346 153176 35402 153232
rect 69662 159296 69718 159352
rect 69570 157936 69626 157992
rect 73434 162016 73490 162072
rect 72882 156576 72938 156632
rect 92386 159296 92442 159352
rect 150530 158752 150586 158808
rect 150438 156032 150494 156088
rect 137098 153992 137154 154048
rect 143354 152904 143410 152960
rect 95146 152496 95202 152552
rect 34242 152360 34298 152416
rect 27526 152224 27582 152280
rect 21362 10920 21418 10976
rect 22098 13096 22154 13152
rect 23110 10240 23166 10296
rect 23754 9424 23810 9480
rect 35990 11600 36046 11656
rect 35898 6840 35954 6896
rect 33874 6160 33930 6216
rect 56506 2352 56562 2408
rect 59174 13640 59230 13696
rect 63590 8200 63646 8256
rect 67638 15816 67694 15872
rect 70674 15816 70730 15872
rect 71778 15136 71834 15192
rect 70674 6024 70730 6080
rect 71042 4800 71098 4856
rect 71778 8064 71834 8120
rect 76102 14728 76158 14784
rect 77206 10784 77262 10840
rect 79230 10648 79286 10704
rect 80150 18672 80206 18728
rect 80150 17312 80206 17368
rect 80610 3712 80666 3768
rect 82082 6568 82138 6624
rect 81346 5072 81402 5128
rect 82450 11736 82506 11792
rect 83186 11600 83242 11656
rect 84382 11872 84438 11928
rect 87142 18672 87198 18728
rect 86958 7928 87014 7984
rect 86682 2488 86738 2544
rect 88430 10240 88486 10296
rect 88430 8880 88486 8936
rect 88338 3984 88394 4040
rect 89534 17176 89590 17232
rect 89534 16360 89590 16416
rect 90730 16224 90786 16280
rect 91374 17992 91430 18048
rect 91098 14864 91154 14920
rect 91190 9288 91246 9344
rect 89810 1128 89866 1184
rect 92570 14592 92626 14648
rect 92570 11600 92626 11656
rect 93122 2080 93178 2136
rect 94134 14864 94190 14920
rect 94594 15136 94650 15192
rect 94410 13776 94466 13832
rect 94962 15272 95018 15328
rect 94962 12280 95018 12336
rect 95146 14728 95202 14784
rect 95146 12416 95202 12472
rect 95238 11872 95294 11928
rect 95238 10240 95294 10296
rect 95790 17176 95846 17232
rect 95790 13504 95846 13560
rect 95790 10784 95846 10840
rect 96342 14728 96398 14784
rect 96342 13640 96398 13696
rect 96526 19216 96582 19272
rect 96526 14456 96582 14512
rect 96526 13640 96582 13696
rect 96526 12960 96582 13016
rect 96526 12144 96582 12200
rect 96250 6704 96306 6760
rect 95238 6160 95294 6216
rect 95054 5344 95110 5400
rect 97354 17720 97410 17776
rect 97170 14592 97226 14648
rect 97078 14456 97134 14512
rect 96894 13776 96950 13832
rect 96802 6568 96858 6624
rect 97814 18128 97870 18184
rect 97814 13504 97870 13560
rect 95238 2760 95294 2816
rect 98182 13232 98238 13288
rect 98090 10920 98146 10976
rect 97998 8064 98054 8120
rect 97998 7520 98054 7576
rect 97998 6840 98054 6896
rect 98734 9424 98790 9480
rect 98458 6568 98514 6624
rect 99470 15272 99526 15328
rect 98826 6432 98882 6488
rect 97630 5480 97686 5536
rect 99562 3304 99618 3360
rect 100298 10512 100354 10568
rect 99746 856 99802 912
rect 100758 17992 100814 18048
rect 100574 15816 100630 15872
rect 100850 12144 100906 12200
rect 101218 15272 101274 15328
rect 101586 16224 101642 16280
rect 101494 11872 101550 11928
rect 100482 5208 100538 5264
rect 101402 8880 101458 8936
rect 100390 1944 100446 2000
rect 93674 176 93730 232
rect 102414 11736 102470 11792
rect 102506 10376 102562 10432
rect 102138 7928 102194 7984
rect 102138 6976 102194 7032
rect 102138 6024 102194 6080
rect 101770 4120 101826 4176
rect 103794 15816 103850 15872
rect 103242 6296 103298 6352
rect 103518 4256 103574 4312
rect 103518 3984 103574 4040
rect 104162 12824 104218 12880
rect 104806 18128 104862 18184
rect 104438 15000 104494 15056
rect 104806 14456 104862 14512
rect 104530 10648 104586 10704
rect 104346 9152 104402 9208
rect 104254 8200 104310 8256
rect 104806 10240 104862 10296
rect 104898 7656 104954 7712
rect 104530 6840 104586 6896
rect 104162 5072 104218 5128
rect 104438 4800 104494 4856
rect 104438 3168 104494 3224
rect 104254 2488 104310 2544
rect 105174 14864 105230 14920
rect 105358 18264 105414 18320
rect 105818 13640 105874 13696
rect 105450 12960 105506 13016
rect 105634 11192 105690 11248
rect 106094 17992 106150 18048
rect 106094 11600 106150 11656
rect 106094 9696 106150 9752
rect 106002 8064 106058 8120
rect 107382 16632 107438 16688
rect 107106 16088 107162 16144
rect 106554 7928 106610 7984
rect 106186 3576 106242 3632
rect 105266 992 105322 1048
rect 107566 15136 107622 15192
rect 107566 13368 107622 13424
rect 107566 13096 107622 13152
rect 107474 12008 107530 12064
rect 107566 11872 107622 11928
rect 107382 10784 107438 10840
rect 107566 6976 107622 7032
rect 107750 18128 107806 18184
rect 108118 16768 108174 16824
rect 107750 12280 107806 12336
rect 108026 7248 108082 7304
rect 107658 6160 107714 6216
rect 108210 5072 108266 5128
rect 108026 4256 108082 4312
rect 107658 2488 107714 2544
rect 108578 11736 108634 11792
rect 109038 10240 109094 10296
rect 108394 6840 108450 6896
rect 110326 16768 110382 16824
rect 109958 15544 110014 15600
rect 110326 15272 110382 15328
rect 110510 18128 110566 18184
rect 110418 11600 110474 11656
rect 110510 11192 110566 11248
rect 110602 9560 110658 9616
rect 110510 8336 110566 8392
rect 110602 6024 110658 6080
rect 111154 15000 111210 15056
rect 111522 18128 111578 18184
rect 111614 17992 111670 18048
rect 111614 17312 111670 17368
rect 111430 14728 111486 14784
rect 111154 12280 111210 12336
rect 111614 11056 111670 11112
rect 109038 3304 109094 3360
rect 109038 2624 109094 2680
rect 110694 3440 110750 3496
rect 110418 2216 110474 2272
rect 111982 9424 112038 9480
rect 111706 3304 111762 3360
rect 111798 3168 111854 3224
rect 111798 1264 111854 1320
rect 113086 18808 113142 18864
rect 112626 11328 112682 11384
rect 113638 18400 113694 18456
rect 113546 16904 113602 16960
rect 113822 14456 113878 14512
rect 113362 9560 113418 9616
rect 113178 9016 113234 9072
rect 113178 8336 113234 8392
rect 113178 5888 113234 5944
rect 112626 2760 112682 2816
rect 114190 17448 114246 17504
rect 114374 13640 114430 13696
rect 114190 12824 114246 12880
rect 114098 11464 114154 11520
rect 114466 13504 114522 13560
rect 114466 12280 114522 12336
rect 114374 9288 114430 9344
rect 114466 7248 114522 7304
rect 114742 17856 114798 17912
rect 114926 17176 114982 17232
rect 114742 15272 114798 15328
rect 114742 13504 114798 13560
rect 114650 8200 114706 8256
rect 114834 7656 114890 7712
rect 115754 16360 115810 16416
rect 116122 14048 116178 14104
rect 115938 12416 115994 12472
rect 115754 11328 115810 11384
rect 115754 10920 115810 10976
rect 115570 7792 115626 7848
rect 115846 7520 115902 7576
rect 115294 6840 115350 6896
rect 114466 6024 114522 6080
rect 117042 13776 117098 13832
rect 114098 3848 114154 3904
rect 113362 2216 113418 2272
rect 115846 2624 115902 2680
rect 117410 17856 117466 17912
rect 117410 15272 117466 15328
rect 117226 13504 117282 13560
rect 117594 15408 117650 15464
rect 117502 12960 117558 13016
rect 118054 17992 118110 18048
rect 117594 10784 117650 10840
rect 117134 9288 117190 9344
rect 118330 13640 118386 13696
rect 118238 13504 118294 13560
rect 118514 18536 118570 18592
rect 118698 17720 118754 17776
rect 118790 17584 118846 17640
rect 119066 17448 119122 17504
rect 118974 15000 119030 15056
rect 118790 14048 118846 14104
rect 118606 12416 118662 12472
rect 119250 10920 119306 10976
rect 119618 17856 119674 17912
rect 119802 17856 119858 17912
rect 118698 6860 118754 6896
rect 118698 6840 118700 6860
rect 118700 6840 118752 6860
rect 118752 6840 118754 6860
rect 119986 12144 120042 12200
rect 119894 9696 119950 9752
rect 120170 17720 120226 17776
rect 120078 9560 120134 9616
rect 117962 2488 118018 2544
rect 118146 2488 118202 2544
rect 120998 19216 121054 19272
rect 120538 7656 120594 7712
rect 120814 16632 120870 16688
rect 121320 19760 121376 19816
rect 121090 15952 121146 16008
rect 120814 5888 120870 5944
rect 121366 12688 121422 12744
rect 121274 9424 121330 9480
rect 121550 15408 121606 15464
rect 122102 19624 122158 19680
rect 121826 17992 121882 18048
rect 122010 15136 122066 15192
rect 121642 4936 121698 4992
rect 122378 17584 122434 17640
rect 122378 15272 122434 15328
rect 122838 17584 122894 17640
rect 123022 18536 123078 18592
rect 122930 16768 122986 16824
rect 123114 17856 123170 17912
rect 123022 15272 123078 15328
rect 123482 17856 123538 17912
rect 122838 13368 122894 13424
rect 123574 16632 123630 16688
rect 122378 3848 122434 3904
rect 122102 2352 122158 2408
rect 122838 1264 122894 1320
rect 123666 13776 123722 13832
rect 124218 17856 124274 17912
rect 125138 18400 125194 18456
rect 125046 17856 125102 17912
rect 124862 17720 124918 17776
rect 124402 15136 124458 15192
rect 124218 13912 124274 13968
rect 124218 13776 124274 13832
rect 124126 11056 124182 11112
rect 124218 8880 124274 8936
rect 123574 2352 123630 2408
rect 124126 1536 124182 1592
rect 125690 17856 125746 17912
rect 125506 17448 125562 17504
rect 126242 17720 126298 17776
rect 126242 15000 126298 15056
rect 125322 13368 125378 13424
rect 125874 13776 125930 13832
rect 126242 12008 126298 12064
rect 126702 19624 126758 19680
rect 126886 16496 126942 16552
rect 126886 11464 126942 11520
rect 126886 10920 126942 10976
rect 127254 19488 127310 19544
rect 127622 17856 127678 17912
rect 127346 17584 127402 17640
rect 127898 19216 127954 19272
rect 127990 18536 128046 18592
rect 128358 18536 128414 18592
rect 128266 16768 128322 16824
rect 127714 7520 127770 7576
rect 128726 17720 128782 17776
rect 128910 17856 128966 17912
rect 129278 17856 129334 17912
rect 128818 16360 128874 16416
rect 129462 17584 129518 17640
rect 129646 18944 129702 19000
rect 129738 16496 129794 16552
rect 129830 15680 129886 15736
rect 129002 13776 129058 13832
rect 128910 10784 128966 10840
rect 127070 2624 127126 2680
rect 126978 1536 127034 1592
rect 126426 40 126482 96
rect 130014 17720 130070 17776
rect 130198 17312 130254 17368
rect 142618 19216 142674 19272
rect 137282 18944 137338 19000
rect 130658 17856 130714 17912
rect 130566 17720 130622 17776
rect 130382 17176 130438 17232
rect 129922 4800 129978 4856
rect 129002 4664 129058 4720
rect 129646 1284 129702 1320
rect 129646 1264 129648 1284
rect 129648 1264 129700 1284
rect 129700 1264 129702 1284
rect 131118 16496 131174 16552
rect 131118 15680 131174 15736
rect 130658 5616 130714 5672
rect 132590 13640 132646 13696
rect 133234 10920 133290 10976
rect 143446 18128 143502 18184
rect 142250 17584 142306 17640
rect 146206 17584 146262 17640
rect 143538 17448 143594 17504
rect 137282 13640 137338 13696
rect 135074 992 135130 1048
rect 136546 1264 136602 1320
rect 140778 8744 140834 8800
rect 140686 6024 140742 6080
rect 143538 5616 143594 5672
rect 145010 2352 145066 2408
rect 147678 17856 147734 17912
rect 150530 13504 150586 13560
rect 149058 11328 149114 11384
rect 147034 6024 147090 6080
rect 146942 4664 146998 4720
rect 146574 2488 146630 2544
rect 150438 3984 150494 4040
rect 151082 155216 151138 155272
rect 150898 151816 150954 151872
rect 151266 153312 151322 153368
rect 150990 19624 151046 19680
rect 150898 12144 150954 12200
rect 151174 9424 151230 9480
rect 152094 153176 152150 153232
rect 152554 153720 152610 153776
rect 153934 153856 153990 153912
rect 157982 153448 158038 153504
rect 156694 152360 156750 152416
rect 160742 152224 160798 152280
rect 152646 16496 152702 16552
rect 153014 17856 153070 17912
rect 153290 19216 153346 19272
rect 153106 17584 153162 17640
rect 153750 15544 153806 15600
rect 152554 9560 152610 9616
rect 154026 18808 154082 18864
rect 153934 16768 153990 16824
rect 154118 11464 154174 11520
rect 154394 15136 154450 15192
rect 154302 13368 154358 13424
rect 154118 8744 154174 8800
rect 155682 16360 155738 16416
rect 155498 13640 155554 13696
rect 155958 12008 156014 12064
rect 157338 12688 157394 12744
rect 156694 10920 156750 10976
rect 169758 159296 169814 159352
rect 163502 157392 163558 157448
rect 162122 153584 162178 153640
rect 160190 3712 160246 3768
rect 209778 151272 209834 151328
rect 240506 16224 240562 16280
rect 253938 16088 253994 16144
rect 299386 19488 299442 19544
rect 302238 18672 302294 18728
rect 298466 14864 298522 14920
rect 299662 2080 299718 2136
rect 306378 18264 306434 18320
rect 313278 1128 313334 1184
rect 329194 5480 329250 5536
rect 335082 1944 335138 2000
rect 340970 5344 341026 5400
rect 371882 160112 371938 160168
rect 345386 176 345442 232
rect 355966 15952 356022 16008
rect 358726 14728 358782 14784
rect 353022 8200 353078 8256
rect 358818 6704 358874 6760
rect 367650 14592 367706 14648
rect 371238 13232 371294 13288
rect 372618 6568 372674 6624
rect 377954 11872 378010 11928
rect 377402 10512 377458 10568
rect 378874 6432 378930 6488
rect 385314 10376 385370 10432
rect 384394 856 384450 912
rect 389454 5208 389510 5264
rect 442262 155080 442318 155136
rect 439502 154128 439558 154184
rect 406566 17312 406622 17368
rect 404266 11736 404322 11792
rect 403714 9288 403770 9344
rect 407210 6296 407266 6352
rect 410798 15816 410854 15872
rect 420918 13096 420974 13152
rect 414294 9152 414350 9208
rect 430578 14456 430634 14512
rect 424966 8064 425022 8120
rect 428462 7928 428518 7984
rect 426162 3576 426218 3632
rect 435546 6160 435602 6216
rect 439134 5072 439190 5128
rect 442630 10240 442686 10296
rect 453210 11600 453266 11656
rect 454498 3440 454554 3496
rect 527178 162016 527234 162072
rect 507858 154944 507914 155000
rect 462318 9016 462374 9072
rect 461582 3304 461638 3360
rect 482374 12960 482430 13016
rect 486422 7792 486478 7848
rect 512642 154808 512698 154864
rect 527178 19352 527234 19408
rect 518346 7656 518402 7712
rect 525430 4936 525486 4992
rect 539598 154672 539654 154728
rect 543738 152088 543794 152144
rect 545118 18536 545174 18592
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580262 670656 580318 670712
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 579894 431568 579950 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245520 580226 245576
rect 579802 232328 579858 232384
rect 579894 219000 579950 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580262 157936 580318 157992
rect 558918 156576 558974 156632
rect 576122 154536 576178 154592
rect 538402 8880 538458 8936
rect 552570 2624 552626 2680
rect 556342 40 556398 96
rect 562322 7520 562378 7576
rect 580262 152632 580318 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 582378 24928 582434 24984
rect 580262 19760 580318 19816
rect 581090 17176 581146 17232
rect 578882 6568 578938 6624
rect 578606 4800 578662 4856
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 73429 162074 73495 162077
rect 527173 162074 527239 162077
rect 73429 162072 527239 162074
rect 73429 162016 73434 162072
rect 73490 162016 527178 162072
rect 527234 162016 527239 162072
rect 73429 162014 527239 162016
rect 73429 162011 73495 162014
rect 527173 162011 527239 162014
rect 9121 160170 9187 160173
rect 371877 160170 371943 160173
rect 9121 160168 371943 160170
rect 9121 160112 9126 160168
rect 9182 160112 371882 160168
rect 371938 160112 371943 160168
rect 9121 160110 371943 160112
rect 9121 160107 9187 160110
rect 371877 160107 371943 160110
rect 18045 159354 18111 159357
rect 69657 159354 69723 159357
rect 18045 159352 69723 159354
rect 18045 159296 18050 159352
rect 18106 159296 69662 159352
rect 69718 159296 69723 159352
rect 18045 159294 69723 159296
rect 18045 159291 18111 159294
rect 69657 159291 69723 159294
rect 92381 159354 92447 159357
rect 169753 159354 169819 159357
rect 92381 159352 169819 159354
rect 92381 159296 92386 159352
rect 92442 159296 169758 159352
rect 169814 159296 169819 159352
rect 92381 159294 169819 159296
rect 92381 159291 92447 159294
rect 169753 159291 169819 159294
rect 20621 158810 20687 158813
rect 150525 158810 150591 158813
rect 20621 158808 150591 158810
rect 20621 158752 20626 158808
rect 20682 158752 150530 158808
rect 150586 158752 150591 158808
rect 20621 158750 150591 158752
rect 20621 158747 20687 158750
rect 150525 158747 150591 158750
rect 69565 157994 69631 157997
rect 580257 157994 580323 157997
rect 69565 157992 580323 157994
rect 69565 157936 69570 157992
rect 69626 157936 580262 157992
rect 580318 157936 580323 157992
rect 69565 157934 580323 157936
rect 69565 157931 69631 157934
rect 580257 157931 580323 157934
rect 18229 157450 18295 157453
rect 163497 157450 163563 157453
rect 18229 157448 163563 157450
rect 18229 157392 18234 157448
rect 18290 157392 163502 157448
rect 163558 157392 163563 157448
rect 18229 157390 163563 157392
rect 18229 157387 18295 157390
rect 163497 157387 163563 157390
rect 72877 156634 72943 156637
rect 558913 156634 558979 156637
rect 72877 156632 558979 156634
rect 72877 156576 72882 156632
rect 72938 156576 558918 156632
rect 558974 156576 558979 156632
rect 72877 156574 558979 156576
rect 72877 156571 72943 156574
rect 558913 156571 558979 156574
rect 14457 156090 14523 156093
rect 150433 156090 150499 156093
rect 14457 156088 150499 156090
rect 14457 156032 14462 156088
rect 14518 156032 150438 156088
rect 150494 156032 150499 156088
rect 14457 156030 150499 156032
rect 14457 156027 14523 156030
rect 150433 156027 150499 156030
rect 22093 155410 22159 155413
rect 35617 155410 35683 155413
rect 22093 155408 35683 155410
rect 22093 155352 22098 155408
rect 22154 155352 35622 155408
rect 35678 155352 35683 155408
rect 22093 155350 35683 155352
rect 22093 155347 22159 155350
rect 35617 155347 35683 155350
rect 31661 155274 31727 155277
rect 151077 155274 151143 155277
rect 31661 155272 151143 155274
rect 31661 155216 31666 155272
rect 31722 155216 151082 155272
rect 151138 155216 151143 155272
rect 31661 155214 151143 155216
rect 31661 155211 31727 155214
rect 151077 155211 151143 155214
rect 19701 155138 19767 155141
rect 442257 155138 442323 155141
rect 19701 155136 442323 155138
rect 19701 155080 19706 155136
rect 19762 155080 442262 155136
rect 442318 155080 442323 155136
rect 19701 155078 442323 155080
rect 19701 155075 19767 155078
rect 442257 155075 442323 155078
rect 19149 155002 19215 155005
rect 507853 155002 507919 155005
rect 19149 155000 507919 155002
rect 19149 154944 19154 155000
rect 19210 154944 507858 155000
rect 507914 154944 507919 155000
rect 19149 154942 507919 154944
rect 19149 154939 19215 154942
rect 507853 154939 507919 154942
rect 19793 154866 19859 154869
rect 512637 154866 512703 154869
rect 19793 154864 512703 154866
rect 19793 154808 19798 154864
rect 19854 154808 512642 154864
rect 512698 154808 512703 154864
rect 19793 154806 512703 154808
rect 19793 154803 19859 154806
rect 512637 154803 512703 154806
rect 14825 154730 14891 154733
rect 539593 154730 539659 154733
rect 14825 154728 539659 154730
rect 14825 154672 14830 154728
rect 14886 154672 539598 154728
rect 539654 154672 539659 154728
rect 14825 154670 539659 154672
rect 14825 154667 14891 154670
rect 539593 154667 539659 154670
rect 28717 154594 28783 154597
rect 576117 154594 576183 154597
rect 28717 154592 576183 154594
rect 28717 154536 28722 154592
rect 28778 154536 576122 154592
rect 576178 154536 576183 154592
rect 28717 154534 576183 154536
rect 28717 154531 28783 154534
rect 576117 154531 576183 154534
rect 28901 154458 28967 154461
rect 31886 154458 31892 154460
rect 28901 154456 31892 154458
rect 28901 154400 28906 154456
rect 28962 154400 31892 154456
rect 28901 154398 31892 154400
rect 28901 154395 28967 154398
rect 31886 154396 31892 154398
rect 31956 154396 31962 154460
rect 14733 154186 14799 154189
rect 439497 154186 439563 154189
rect 14733 154184 439563 154186
rect 14733 154128 14738 154184
rect 14794 154128 439502 154184
rect 439558 154128 439563 154184
rect 14733 154126 439563 154128
rect 14733 154123 14799 154126
rect 439497 154123 439563 154126
rect 34973 154050 35039 154053
rect 137093 154050 137159 154053
rect 34973 154048 137159 154050
rect 34973 153992 34978 154048
rect 35034 153992 137098 154048
rect 137154 153992 137159 154048
rect 34973 153990 137159 153992
rect 34973 153987 35039 153990
rect 137093 153987 137159 153990
rect 29821 153914 29887 153917
rect 153929 153914 153995 153917
rect 29821 153912 153995 153914
rect 29821 153856 29826 153912
rect 29882 153856 153934 153912
rect 153990 153856 153995 153912
rect 29821 153854 153995 153856
rect 29821 153851 29887 153854
rect 153929 153851 153995 153854
rect 13629 153778 13695 153781
rect 22093 153778 22159 153781
rect 13629 153776 22159 153778
rect 13629 153720 13634 153776
rect 13690 153720 22098 153776
rect 22154 153720 22159 153776
rect 13629 153718 22159 153720
rect 13629 153715 13695 153718
rect 22093 153715 22159 153718
rect 26141 153778 26207 153781
rect 152549 153778 152615 153781
rect 26141 153776 152615 153778
rect 26141 153720 26146 153776
rect 26202 153720 152554 153776
rect 152610 153720 152615 153776
rect 26141 153718 152615 153720
rect 26141 153715 26207 153718
rect 152549 153715 152615 153718
rect 22185 153642 22251 153645
rect 25814 153642 25820 153644
rect 22185 153640 25820 153642
rect 22185 153584 22190 153640
rect 22246 153584 25820 153640
rect 22185 153582 25820 153584
rect 22185 153579 22251 153582
rect 25814 153580 25820 153582
rect 25884 153580 25890 153644
rect 30833 153642 30899 153645
rect 162117 153642 162183 153645
rect 30833 153640 162183 153642
rect 30833 153584 30838 153640
rect 30894 153584 162122 153640
rect 162178 153584 162183 153640
rect 30833 153582 162183 153584
rect 30833 153579 30899 153582
rect 162117 153579 162183 153582
rect 24301 153506 24367 153509
rect 157977 153506 158043 153509
rect 24301 153504 158043 153506
rect 24301 153448 24306 153504
rect 24362 153448 157982 153504
rect 158038 153448 158043 153504
rect 24301 153446 158043 153448
rect 24301 153443 24367 153446
rect 157977 153443 158043 153446
rect 14549 153370 14615 153373
rect 151261 153370 151327 153373
rect 14549 153368 151327 153370
rect 14549 153312 14554 153368
rect 14610 153312 151266 153368
rect 151322 153312 151327 153368
rect 14549 153310 151327 153312
rect 14549 153307 14615 153310
rect 151261 153307 151327 153310
rect 13537 153234 13603 153237
rect 35341 153234 35407 153237
rect 13537 153232 35407 153234
rect 13537 153176 13542 153232
rect 13598 153176 35346 153232
rect 35402 153176 35407 153232
rect 13537 153174 35407 153176
rect 13537 153171 13603 153174
rect 35341 153171 35407 153174
rect 143574 153172 143580 153236
rect 143644 153234 143650 153236
rect 152089 153234 152155 153237
rect 143644 153232 152155 153234
rect 143644 153176 152094 153232
rect 152150 153176 152155 153232
rect 143644 153174 152155 153176
rect 143644 153172 143650 153174
rect 152089 153171 152155 153174
rect 139342 152900 139348 152964
rect 139412 152962 139418 152964
rect 143349 152962 143415 152965
rect 139412 152960 143415 152962
rect 139412 152904 143354 152960
rect 143410 152904 143415 152960
rect 139412 152902 143415 152904
rect 139412 152900 139418 152902
rect 143349 152899 143415 152902
rect 25405 152690 25471 152693
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 25405 152688 580323 152690
rect 25405 152632 25410 152688
rect 25466 152632 580262 152688
rect 580318 152632 580323 152688
rect 25405 152630 580323 152632
rect 25405 152627 25471 152630
rect 580257 152627 580323 152630
rect 583342 152630 584960 152690
rect 33041 152554 33107 152557
rect 95141 152554 95207 152557
rect 137870 152554 137876 152556
rect 33041 152552 45570 152554
rect 33041 152496 33046 152552
rect 33102 152496 45570 152552
rect 33041 152494 45570 152496
rect 33041 152491 33107 152494
rect 34237 152418 34303 152421
rect 37590 152418 37596 152420
rect 34237 152416 37596 152418
rect 34237 152360 34242 152416
rect 34298 152360 37596 152416
rect 34237 152358 37596 152360
rect 34237 152355 34303 152358
rect 37590 152356 37596 152358
rect 37660 152356 37666 152420
rect 45510 152418 45570 152494
rect 95141 152552 137876 152554
rect 95141 152496 95146 152552
rect 95202 152496 137876 152552
rect 95141 152494 137876 152496
rect 95141 152491 95207 152494
rect 137870 152492 137876 152494
rect 137940 152492 137946 152556
rect 583342 152554 583402 152630
rect 583520 152554 584960 152630
rect 583342 152540 584960 152554
rect 583342 152494 583586 152540
rect 156689 152418 156755 152421
rect 45510 152416 156755 152418
rect 45510 152360 156694 152416
rect 156750 152360 156755 152416
rect 45510 152358 156755 152360
rect 156689 152355 156755 152358
rect 27521 152282 27587 152285
rect 160737 152282 160803 152285
rect 27521 152280 160803 152282
rect 27521 152224 27526 152280
rect 27582 152224 160742 152280
rect 160798 152224 160803 152280
rect 27521 152222 160803 152224
rect 27521 152219 27587 152222
rect 160737 152219 160803 152222
rect 19926 152084 19932 152148
rect 19996 152146 20002 152148
rect 543733 152146 543799 152149
rect 19996 152144 543799 152146
rect 19996 152088 543738 152144
rect 543794 152088 543799 152144
rect 19996 152086 543799 152088
rect 19996 152084 20002 152086
rect 543733 152083 543799 152086
rect 37590 151948 37596 152012
rect 37660 152010 37666 152012
rect 583526 152010 583586 152494
rect 37660 151950 583586 152010
rect 37660 151948 37666 151950
rect 10501 151874 10567 151877
rect 35750 151874 35756 151876
rect 10501 151872 35756 151874
rect 10501 151816 10506 151872
rect 10562 151816 35756 151872
rect 10501 151814 35756 151816
rect 10501 151811 10567 151814
rect 35750 151812 35756 151814
rect 35820 151812 35826 151876
rect 136582 151812 136588 151876
rect 136652 151874 136658 151876
rect 150893 151874 150959 151877
rect 136652 151872 150959 151874
rect 136652 151816 150898 151872
rect 150954 151816 150959 151872
rect 136652 151814 150959 151816
rect 136652 151812 136658 151814
rect 150893 151811 150959 151814
rect 25814 151676 25820 151740
rect 25884 151738 25890 151740
rect 143574 151738 143580 151740
rect 25884 151678 143580 151738
rect 25884 151676 25890 151678
rect 143574 151676 143580 151678
rect 143644 151676 143650 151740
rect 31886 151540 31892 151604
rect 31956 151602 31962 151604
rect 136582 151602 136588 151604
rect 31956 151542 136588 151602
rect 31956 151540 31962 151542
rect 136582 151540 136588 151542
rect 136652 151540 136658 151604
rect 35750 151404 35756 151468
rect 35820 151466 35826 151468
rect 139342 151466 139348 151468
rect 35820 151406 139348 151466
rect 35820 151404 35826 151406
rect 139342 151404 139348 151406
rect 139412 151404 139418 151468
rect 137870 151268 137876 151332
rect 137940 151330 137946 151332
rect 209773 151330 209839 151333
rect 137940 151328 209839 151330
rect 137940 151272 209778 151328
rect 209834 151272 209839 151328
rect 137940 151270 209839 151272
rect 137940 151268 137946 151270
rect 209773 151267 209839 151270
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3141 97610 3207 97613
rect -960 97608 3207 97610
rect -960 97552 3146 97608
rect 3202 97552 3207 97608
rect -960 97550 3207 97552
rect -960 97460 480 97550
rect 3141 97547 3207 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2957 84690 3023 84693
rect -960 84688 3023 84690
rect -960 84632 2962 84688
rect 3018 84632 3023 84688
rect -960 84630 3023 84632
rect -960 84540 480 84630
rect 2957 84627 3023 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 151118 24924 151124 24988
rect 151188 24986 151194 24988
rect 582373 24986 582439 24989
rect 151188 24984 582439 24986
rect 151188 24928 582378 24984
rect 582434 24928 582439 24984
rect 151188 24926 582439 24928
rect 151188 24924 151194 24926
rect 582373 24923 582439 24926
rect 16021 19954 16087 19957
rect 16021 19952 103530 19954
rect 16021 19896 16026 19952
rect 16082 19896 103530 19952
rect 16021 19894 103530 19896
rect 16021 19891 16087 19894
rect 103470 19818 103530 19894
rect 121315 19818 121381 19821
rect 103470 19816 121381 19818
rect 103470 19760 121320 19816
rect 121376 19760 121381 19816
rect 103470 19758 121381 19760
rect 121315 19755 121381 19758
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 122097 19682 122163 19685
rect 126697 19682 126763 19685
rect 150985 19682 151051 19685
rect 122097 19680 122850 19682
rect 122097 19624 122102 19680
rect 122158 19624 122850 19680
rect 122097 19622 122850 19624
rect 122097 19619 122163 19622
rect -960 19410 480 19500
rect 3141 19410 3207 19413
rect -960 19408 3207 19410
rect -960 19352 3146 19408
rect 3202 19352 3207 19408
rect -960 19350 3207 19352
rect 122790 19410 122850 19622
rect 126697 19680 151051 19682
rect 126697 19624 126702 19680
rect 126758 19624 150990 19680
rect 151046 19624 151051 19680
rect 583520 19668 584960 19758
rect 126697 19622 151051 19624
rect 126697 19619 126763 19622
rect 150985 19619 151051 19622
rect 127249 19546 127315 19549
rect 299381 19546 299447 19549
rect 127249 19544 299447 19546
rect 127249 19488 127254 19544
rect 127310 19488 299386 19544
rect 299442 19488 299447 19544
rect 127249 19486 299447 19488
rect 127249 19483 127315 19486
rect 299381 19483 299447 19486
rect 527173 19410 527239 19413
rect 122790 19408 527239 19410
rect 122790 19352 527178 19408
rect 527234 19352 527239 19408
rect 122790 19350 527239 19352
rect -960 19260 480 19350
rect 3141 19347 3207 19350
rect 527173 19347 527239 19350
rect 19701 19274 19767 19277
rect 96521 19274 96587 19277
rect 19701 19272 96587 19274
rect 19701 19216 19706 19272
rect 19762 19216 96526 19272
rect 96582 19216 96587 19272
rect 19701 19214 96587 19216
rect 19701 19211 19767 19214
rect 96521 19211 96587 19214
rect 120993 19274 121059 19277
rect 127893 19274 127959 19277
rect 120993 19272 127959 19274
rect 120993 19216 120998 19272
rect 121054 19216 127898 19272
rect 127954 19216 127959 19272
rect 120993 19214 127959 19216
rect 120993 19211 121059 19214
rect 127893 19211 127959 19214
rect 142613 19274 142679 19277
rect 153285 19274 153351 19277
rect 142613 19272 153351 19274
rect 142613 19216 142618 19272
rect 142674 19216 153290 19272
rect 153346 19216 153351 19272
rect 142613 19214 153351 19216
rect 142613 19211 142679 19214
rect 153285 19211 153351 19214
rect 129641 19002 129707 19005
rect 137277 19002 137343 19005
rect 129641 19000 137343 19002
rect 129641 18944 129646 19000
rect 129702 18944 137282 19000
rect 137338 18944 137343 19000
rect 129641 18942 137343 18944
rect 129641 18939 129707 18942
rect 137277 18939 137343 18942
rect 113081 18866 113147 18869
rect 154021 18866 154087 18869
rect 113081 18864 154087 18866
rect 113081 18808 113086 18864
rect 113142 18808 154026 18864
rect 154082 18808 154087 18864
rect 113081 18806 154087 18808
rect 113081 18803 113147 18806
rect 154021 18803 154087 18806
rect 17677 18730 17743 18733
rect 80145 18730 80211 18733
rect 17677 18728 80211 18730
rect 17677 18672 17682 18728
rect 17738 18672 80150 18728
rect 80206 18672 80211 18728
rect 17677 18670 80211 18672
rect 17677 18667 17743 18670
rect 80145 18667 80211 18670
rect 87137 18730 87203 18733
rect 302233 18730 302299 18733
rect 87137 18728 302299 18730
rect 87137 18672 87142 18728
rect 87198 18672 302238 18728
rect 302294 18672 302299 18728
rect 87137 18670 302299 18672
rect 87137 18667 87203 18670
rect 302233 18667 302299 18670
rect 17401 18594 17467 18597
rect 118509 18594 118575 18597
rect 17401 18592 118575 18594
rect 17401 18536 17406 18592
rect 17462 18536 118514 18592
rect 118570 18536 118575 18592
rect 17401 18534 118575 18536
rect 17401 18531 17467 18534
rect 118509 18531 118575 18534
rect 123017 18594 123083 18597
rect 127985 18594 128051 18597
rect 123017 18592 128051 18594
rect 123017 18536 123022 18592
rect 123078 18536 127990 18592
rect 128046 18536 128051 18592
rect 123017 18534 128051 18536
rect 123017 18531 123083 18534
rect 127985 18531 128051 18534
rect 128353 18594 128419 18597
rect 545113 18594 545179 18597
rect 128353 18592 545179 18594
rect 128353 18536 128358 18592
rect 128414 18536 545118 18592
rect 545174 18536 545179 18592
rect 128353 18534 545179 18536
rect 128353 18531 128419 18534
rect 545113 18531 545179 18534
rect 113633 18458 113699 18461
rect 125133 18458 125199 18461
rect 113633 18456 125199 18458
rect 113633 18400 113638 18456
rect 113694 18400 125138 18456
rect 125194 18400 125199 18456
rect 113633 18398 125199 18400
rect 113633 18395 113699 18398
rect 125133 18395 125199 18398
rect 105353 18322 105419 18325
rect 306373 18322 306439 18325
rect 105353 18320 306439 18322
rect 105353 18264 105358 18320
rect 105414 18264 306378 18320
rect 306434 18264 306439 18320
rect 105353 18262 306439 18264
rect 105353 18259 105419 18262
rect 306373 18259 306439 18262
rect 97809 18186 97875 18189
rect 104801 18186 104867 18189
rect 97809 18184 104867 18186
rect 97809 18128 97814 18184
rect 97870 18128 104806 18184
rect 104862 18128 104867 18184
rect 97809 18126 104867 18128
rect 97809 18123 97875 18126
rect 104801 18123 104867 18126
rect 107745 18186 107811 18189
rect 110505 18186 110571 18189
rect 107745 18184 110571 18186
rect 107745 18128 107750 18184
rect 107806 18128 110510 18184
rect 110566 18128 110571 18184
rect 107745 18126 110571 18128
rect 107745 18123 107811 18126
rect 110505 18123 110571 18126
rect 111517 18186 111583 18189
rect 143441 18186 143507 18189
rect 111517 18184 143507 18186
rect 111517 18128 111522 18184
rect 111578 18128 143446 18184
rect 143502 18128 143507 18184
rect 111517 18126 143507 18128
rect 111517 18123 111583 18126
rect 143441 18123 143507 18126
rect 91369 18050 91435 18053
rect 100753 18050 100819 18053
rect 91369 18048 100819 18050
rect 91369 17992 91374 18048
rect 91430 17992 100758 18048
rect 100814 17992 100819 18048
rect 91369 17990 100819 17992
rect 91369 17987 91435 17990
rect 100753 17987 100819 17990
rect 106089 18050 106155 18053
rect 111609 18050 111675 18053
rect 106089 18048 111675 18050
rect 106089 17992 106094 18048
rect 106150 17992 111614 18048
rect 111670 17992 111675 18048
rect 106089 17990 111675 17992
rect 106089 17987 106155 17990
rect 111609 17987 111675 17990
rect 118049 18050 118115 18053
rect 121821 18050 121887 18053
rect 118049 18048 121887 18050
rect 118049 17992 118054 18048
rect 118110 17992 121826 18048
rect 121882 17992 121887 18048
rect 118049 17990 121887 17992
rect 118049 17987 118115 17990
rect 121821 17987 121887 17990
rect 18873 17914 18939 17917
rect 114737 17914 114803 17917
rect 18873 17912 114803 17914
rect 18873 17856 18878 17912
rect 18934 17856 114742 17912
rect 114798 17856 114803 17912
rect 18873 17854 114803 17856
rect 18873 17851 18939 17854
rect 114737 17851 114803 17854
rect 117405 17914 117471 17917
rect 119613 17914 119679 17917
rect 117405 17912 119679 17914
rect 117405 17856 117410 17912
rect 117466 17856 119618 17912
rect 119674 17856 119679 17912
rect 117405 17854 119679 17856
rect 117405 17851 117471 17854
rect 119613 17851 119679 17854
rect 119797 17914 119863 17917
rect 123109 17914 123175 17917
rect 119797 17912 123175 17914
rect 119797 17856 119802 17912
rect 119858 17856 123114 17912
rect 123170 17856 123175 17912
rect 119797 17854 123175 17856
rect 119797 17851 119863 17854
rect 123109 17851 123175 17854
rect 123477 17914 123543 17917
rect 124213 17914 124279 17917
rect 123477 17912 124279 17914
rect 123477 17856 123482 17912
rect 123538 17856 124218 17912
rect 124274 17856 124279 17912
rect 123477 17854 124279 17856
rect 123477 17851 123543 17854
rect 124213 17851 124279 17854
rect 125041 17914 125107 17917
rect 125685 17914 125751 17917
rect 125041 17912 125751 17914
rect 125041 17856 125046 17912
rect 125102 17856 125690 17912
rect 125746 17856 125751 17912
rect 125041 17854 125751 17856
rect 125041 17851 125107 17854
rect 125685 17851 125751 17854
rect 127617 17914 127683 17917
rect 128905 17914 128971 17917
rect 127617 17912 128971 17914
rect 127617 17856 127622 17912
rect 127678 17856 128910 17912
rect 128966 17856 128971 17912
rect 127617 17854 128971 17856
rect 127617 17851 127683 17854
rect 128905 17851 128971 17854
rect 129273 17914 129339 17917
rect 130653 17914 130719 17917
rect 129273 17912 130719 17914
rect 129273 17856 129278 17912
rect 129334 17856 130658 17912
rect 130714 17856 130719 17912
rect 129273 17854 130719 17856
rect 129273 17851 129339 17854
rect 130653 17851 130719 17854
rect 147673 17914 147739 17917
rect 153009 17914 153075 17917
rect 147673 17912 153075 17914
rect 147673 17856 147678 17912
rect 147734 17856 153014 17912
rect 153070 17856 153075 17912
rect 147673 17854 153075 17856
rect 147673 17851 147739 17854
rect 153009 17851 153075 17854
rect 17677 17778 17743 17781
rect 97349 17778 97415 17781
rect 17677 17776 97415 17778
rect 17677 17720 17682 17776
rect 17738 17720 97354 17776
rect 97410 17720 97415 17776
rect 17677 17718 97415 17720
rect 17677 17715 17743 17718
rect 97349 17715 97415 17718
rect 118693 17778 118759 17781
rect 120165 17778 120231 17781
rect 118693 17776 120231 17778
rect 118693 17720 118698 17776
rect 118754 17720 120170 17776
rect 120226 17720 120231 17776
rect 118693 17718 120231 17720
rect 118693 17715 118759 17718
rect 120165 17715 120231 17718
rect 124857 17778 124923 17781
rect 126237 17778 126303 17781
rect 124857 17776 126303 17778
rect 124857 17720 124862 17776
rect 124918 17720 126242 17776
rect 126298 17720 126303 17776
rect 124857 17718 126303 17720
rect 124857 17715 124923 17718
rect 126237 17715 126303 17718
rect 128721 17778 128787 17781
rect 130009 17778 130075 17781
rect 128721 17776 130075 17778
rect 128721 17720 128726 17776
rect 128782 17720 130014 17776
rect 130070 17720 130075 17776
rect 128721 17718 130075 17720
rect 128721 17715 128787 17718
rect 130009 17715 130075 17718
rect 130561 17778 130627 17781
rect 151118 17778 151124 17780
rect 130561 17776 151124 17778
rect 130561 17720 130566 17776
rect 130622 17720 151124 17776
rect 130561 17718 151124 17720
rect 130561 17715 130627 17718
rect 151118 17716 151124 17718
rect 151188 17716 151194 17780
rect 118785 17642 118851 17645
rect 122373 17642 122439 17645
rect 118785 17640 122439 17642
rect 118785 17584 118790 17640
rect 118846 17584 122378 17640
rect 122434 17584 122439 17640
rect 118785 17582 122439 17584
rect 118785 17579 118851 17582
rect 122373 17579 122439 17582
rect 122833 17642 122899 17645
rect 127341 17642 127407 17645
rect 122833 17640 127407 17642
rect 122833 17584 122838 17640
rect 122894 17584 127346 17640
rect 127402 17584 127407 17640
rect 122833 17582 127407 17584
rect 122833 17579 122899 17582
rect 127341 17579 127407 17582
rect 129457 17642 129523 17645
rect 142245 17642 142311 17645
rect 129457 17640 142311 17642
rect 129457 17584 129462 17640
rect 129518 17584 142250 17640
rect 142306 17584 142311 17640
rect 129457 17582 142311 17584
rect 129457 17579 129523 17582
rect 142245 17579 142311 17582
rect 146201 17642 146267 17645
rect 153101 17642 153167 17645
rect 146201 17640 153167 17642
rect 146201 17584 146206 17640
rect 146262 17584 153106 17640
rect 153162 17584 153167 17640
rect 146201 17582 153167 17584
rect 146201 17579 146267 17582
rect 153101 17579 153167 17582
rect 114185 17506 114251 17509
rect 119061 17506 119127 17509
rect 114185 17504 119127 17506
rect 114185 17448 114190 17504
rect 114246 17448 119066 17504
rect 119122 17448 119127 17504
rect 114185 17446 119127 17448
rect 114185 17443 114251 17446
rect 119061 17443 119127 17446
rect 125501 17506 125567 17509
rect 143533 17506 143599 17509
rect 125501 17504 143599 17506
rect 125501 17448 125506 17504
rect 125562 17448 143538 17504
rect 143594 17448 143599 17504
rect 125501 17446 143599 17448
rect 125501 17443 125567 17446
rect 143533 17443 143599 17446
rect 80145 17370 80211 17373
rect 111609 17370 111675 17373
rect 80145 17368 111675 17370
rect 80145 17312 80150 17368
rect 80206 17312 111614 17368
rect 111670 17312 111675 17368
rect 80145 17310 111675 17312
rect 80145 17307 80211 17310
rect 111609 17307 111675 17310
rect 130193 17370 130259 17373
rect 406561 17370 406627 17373
rect 130193 17368 406627 17370
rect 130193 17312 130198 17368
rect 130254 17312 406566 17368
rect 406622 17312 406627 17368
rect 130193 17310 406627 17312
rect 130193 17307 130259 17310
rect 406561 17307 406627 17310
rect 18965 17234 19031 17237
rect 89529 17234 89595 17237
rect 18965 17232 89595 17234
rect 18965 17176 18970 17232
rect 19026 17176 89534 17232
rect 89590 17176 89595 17232
rect 18965 17174 89595 17176
rect 18965 17171 19031 17174
rect 89529 17171 89595 17174
rect 95785 17234 95851 17237
rect 114921 17234 114987 17237
rect 95785 17232 114987 17234
rect 95785 17176 95790 17232
rect 95846 17176 114926 17232
rect 114982 17176 114987 17232
rect 95785 17174 114987 17176
rect 95785 17171 95851 17174
rect 114921 17171 114987 17174
rect 130377 17234 130443 17237
rect 581085 17234 581151 17237
rect 130377 17232 581151 17234
rect 130377 17176 130382 17232
rect 130438 17176 581090 17232
rect 581146 17176 581151 17232
rect 130377 17174 581151 17176
rect 130377 17171 130443 17174
rect 581085 17171 581151 17174
rect 113541 16962 113607 16965
rect 108990 16960 113607 16962
rect 108990 16904 113546 16960
rect 113602 16904 113607 16960
rect 108990 16902 113607 16904
rect 108113 16826 108179 16829
rect 108990 16826 109050 16902
rect 113541 16899 113607 16902
rect 108113 16824 109050 16826
rect 108113 16768 108118 16824
rect 108174 16768 109050 16824
rect 108113 16766 109050 16768
rect 110321 16826 110387 16829
rect 122925 16826 122991 16829
rect 110321 16824 122991 16826
rect 110321 16768 110326 16824
rect 110382 16768 122930 16824
rect 122986 16768 122991 16824
rect 110321 16766 122991 16768
rect 108113 16763 108179 16766
rect 110321 16763 110387 16766
rect 122925 16763 122991 16766
rect 128261 16826 128327 16829
rect 153929 16826 153995 16829
rect 128261 16824 153995 16826
rect 128261 16768 128266 16824
rect 128322 16768 153934 16824
rect 153990 16768 153995 16824
rect 128261 16766 153995 16768
rect 128261 16763 128327 16766
rect 153929 16763 153995 16766
rect 13169 16690 13235 16693
rect 18689 16690 18755 16693
rect 107377 16690 107443 16693
rect 13169 16688 18755 16690
rect 13169 16632 13174 16688
rect 13230 16632 18694 16688
rect 18750 16632 18755 16688
rect 13169 16630 18755 16632
rect 13169 16627 13235 16630
rect 18689 16627 18755 16630
rect 96570 16688 107443 16690
rect 96570 16632 107382 16688
rect 107438 16632 107443 16688
rect 96570 16630 107443 16632
rect 14825 16554 14891 16557
rect 96570 16554 96630 16630
rect 107377 16627 107443 16630
rect 120809 16690 120875 16693
rect 123569 16690 123635 16693
rect 120809 16688 123635 16690
rect 120809 16632 120814 16688
rect 120870 16632 123574 16688
rect 123630 16632 123635 16688
rect 120809 16630 123635 16632
rect 120809 16627 120875 16630
rect 123569 16627 123635 16630
rect 14825 16552 96630 16554
rect 14825 16496 14830 16552
rect 14886 16496 96630 16552
rect 14825 16494 96630 16496
rect 126881 16554 126947 16557
rect 129733 16554 129799 16557
rect 126881 16552 129799 16554
rect 126881 16496 126886 16552
rect 126942 16496 129738 16552
rect 129794 16496 129799 16552
rect 126881 16494 129799 16496
rect 14825 16491 14891 16494
rect 126881 16491 126947 16494
rect 129733 16491 129799 16494
rect 131113 16554 131179 16557
rect 152641 16554 152707 16557
rect 131113 16552 152707 16554
rect 131113 16496 131118 16552
rect 131174 16496 152646 16552
rect 152702 16496 152707 16552
rect 131113 16494 152707 16496
rect 131113 16491 131179 16494
rect 152641 16491 152707 16494
rect 89529 16418 89595 16421
rect 115749 16418 115815 16421
rect 89529 16416 115815 16418
rect 89529 16360 89534 16416
rect 89590 16360 115754 16416
rect 115810 16360 115815 16416
rect 89529 16358 115815 16360
rect 89529 16355 89595 16358
rect 115749 16355 115815 16358
rect 128813 16418 128879 16421
rect 155677 16418 155743 16421
rect 128813 16416 155743 16418
rect 128813 16360 128818 16416
rect 128874 16360 155682 16416
rect 155738 16360 155743 16416
rect 128813 16358 155743 16360
rect 128813 16355 128879 16358
rect 155677 16355 155743 16358
rect 20161 16282 20227 16285
rect 90725 16282 90791 16285
rect 20161 16280 90791 16282
rect 20161 16224 20166 16280
rect 20222 16224 90730 16280
rect 90786 16224 90791 16280
rect 20161 16222 90791 16224
rect 20161 16219 20227 16222
rect 90725 16219 90791 16222
rect 101581 16282 101647 16285
rect 240501 16282 240567 16285
rect 101581 16280 240567 16282
rect 101581 16224 101586 16280
rect 101642 16224 240506 16280
rect 240562 16224 240567 16280
rect 101581 16222 240567 16224
rect 101581 16219 101647 16222
rect 240501 16219 240567 16222
rect 107101 16146 107167 16149
rect 253933 16146 253999 16149
rect 107101 16144 253999 16146
rect 107101 16088 107106 16144
rect 107162 16088 253938 16144
rect 253994 16088 253999 16144
rect 107101 16086 253999 16088
rect 107101 16083 107167 16086
rect 253933 16083 253999 16086
rect 121085 16010 121151 16013
rect 355961 16010 356027 16013
rect 121085 16008 356027 16010
rect 121085 15952 121090 16008
rect 121146 15952 355966 16008
rect 356022 15952 356027 16008
rect 121085 15950 356027 15952
rect 121085 15947 121151 15950
rect 355961 15947 356027 15950
rect 14733 15874 14799 15877
rect 67633 15874 67699 15877
rect 14733 15872 67699 15874
rect 14733 15816 14738 15872
rect 14794 15816 67638 15872
rect 67694 15816 67699 15872
rect 14733 15814 67699 15816
rect 14733 15811 14799 15814
rect 67633 15811 67699 15814
rect 70669 15874 70735 15877
rect 100569 15874 100635 15877
rect 70669 15872 100635 15874
rect 70669 15816 70674 15872
rect 70730 15816 100574 15872
rect 100630 15816 100635 15872
rect 70669 15814 100635 15816
rect 70669 15811 70735 15814
rect 100569 15811 100635 15814
rect 103789 15874 103855 15877
rect 410793 15874 410859 15877
rect 103789 15872 410859 15874
rect 103789 15816 103794 15872
rect 103850 15816 410798 15872
rect 410854 15816 410859 15872
rect 103789 15814 410859 15816
rect 103789 15811 103855 15814
rect 410793 15811 410859 15814
rect 129825 15738 129891 15741
rect 131113 15738 131179 15741
rect 129825 15736 131179 15738
rect 129825 15680 129830 15736
rect 129886 15680 131118 15736
rect 131174 15680 131179 15736
rect 129825 15678 131179 15680
rect 129825 15675 129891 15678
rect 131113 15675 131179 15678
rect 109953 15602 110019 15605
rect 153745 15602 153811 15605
rect 109953 15600 153811 15602
rect 109953 15544 109958 15600
rect 110014 15544 153750 15600
rect 153806 15544 153811 15600
rect 109953 15542 153811 15544
rect 109953 15539 110019 15542
rect 153745 15539 153811 15542
rect 117589 15466 117655 15469
rect 121545 15466 121611 15469
rect 117589 15464 121611 15466
rect 117589 15408 117594 15464
rect 117650 15408 121550 15464
rect 121606 15408 121611 15464
rect 117589 15406 121611 15408
rect 117589 15403 117655 15406
rect 121545 15403 121611 15406
rect 94957 15330 95023 15333
rect 99465 15330 99531 15333
rect 101213 15330 101279 15333
rect 110321 15330 110387 15333
rect 94957 15328 99531 15330
rect 94957 15272 94962 15328
rect 95018 15272 99470 15328
rect 99526 15272 99531 15328
rect 94957 15270 99531 15272
rect 94957 15267 95023 15270
rect 99465 15267 99531 15270
rect 99606 15328 101279 15330
rect 99606 15272 101218 15328
rect 101274 15272 101279 15328
rect 99606 15270 101279 15272
rect 9489 15194 9555 15197
rect 71773 15194 71839 15197
rect 9489 15192 71839 15194
rect 9489 15136 9494 15192
rect 9550 15136 71778 15192
rect 71834 15136 71839 15192
rect 9489 15134 71839 15136
rect 9489 15131 9555 15134
rect 71773 15131 71839 15134
rect 94589 15194 94655 15197
rect 99606 15194 99666 15270
rect 101213 15267 101279 15270
rect 104942 15328 110387 15330
rect 104942 15272 110326 15328
rect 110382 15272 110387 15328
rect 104942 15270 110387 15272
rect 104942 15194 105002 15270
rect 110321 15267 110387 15270
rect 114737 15330 114803 15333
rect 117405 15330 117471 15333
rect 114737 15328 117471 15330
rect 114737 15272 114742 15328
rect 114798 15272 117410 15328
rect 117466 15272 117471 15328
rect 114737 15270 117471 15272
rect 114737 15267 114803 15270
rect 117405 15267 117471 15270
rect 122373 15330 122439 15333
rect 123017 15330 123083 15333
rect 122373 15328 123083 15330
rect 122373 15272 122378 15328
rect 122434 15272 123022 15328
rect 123078 15272 123083 15328
rect 122373 15270 123083 15272
rect 122373 15267 122439 15270
rect 123017 15267 123083 15270
rect 94589 15192 99666 15194
rect 94589 15136 94594 15192
rect 94650 15136 99666 15192
rect 94589 15134 99666 15136
rect 103470 15134 105002 15194
rect 107561 15194 107627 15197
rect 122005 15194 122071 15197
rect 107561 15192 122071 15194
rect 107561 15136 107566 15192
rect 107622 15136 122010 15192
rect 122066 15136 122071 15192
rect 107561 15134 122071 15136
rect 94589 15131 94655 15134
rect 91093 14922 91159 14925
rect 94129 14922 94195 14925
rect 91093 14920 94195 14922
rect 91093 14864 91098 14920
rect 91154 14864 94134 14920
rect 94190 14864 94195 14920
rect 91093 14862 94195 14864
rect 91093 14859 91159 14862
rect 94129 14859 94195 14862
rect 76097 14786 76163 14789
rect 95141 14786 95207 14789
rect 76097 14784 95207 14786
rect 76097 14728 76102 14784
rect 76158 14728 95146 14784
rect 95202 14728 95207 14784
rect 76097 14726 95207 14728
rect 76097 14723 76163 14726
rect 95141 14723 95207 14726
rect 96337 14786 96403 14789
rect 103470 14786 103530 15134
rect 107561 15131 107627 15134
rect 122005 15131 122071 15134
rect 124397 15194 124463 15197
rect 154389 15194 154455 15197
rect 124397 15192 154455 15194
rect 124397 15136 124402 15192
rect 124458 15136 154394 15192
rect 154450 15136 154455 15192
rect 124397 15134 154455 15136
rect 124397 15131 124463 15134
rect 154389 15131 154455 15134
rect 104433 15058 104499 15061
rect 111149 15058 111215 15061
rect 104433 15056 111215 15058
rect 104433 15000 104438 15056
rect 104494 15000 111154 15056
rect 111210 15000 111215 15056
rect 104433 14998 111215 15000
rect 104433 14995 104499 14998
rect 111149 14995 111215 14998
rect 118969 15058 119035 15061
rect 126237 15058 126303 15061
rect 118969 15056 126303 15058
rect 118969 15000 118974 15056
rect 119030 15000 126242 15056
rect 126298 15000 126303 15056
rect 118969 14998 126303 15000
rect 118969 14995 119035 14998
rect 126237 14995 126303 14998
rect 105169 14922 105235 14925
rect 298461 14922 298527 14925
rect 105169 14920 298527 14922
rect 105169 14864 105174 14920
rect 105230 14864 298466 14920
rect 298522 14864 298527 14920
rect 105169 14862 298527 14864
rect 105169 14859 105235 14862
rect 298461 14859 298527 14862
rect 96337 14784 103530 14786
rect 96337 14728 96342 14784
rect 96398 14728 103530 14784
rect 96337 14726 103530 14728
rect 111425 14786 111491 14789
rect 358721 14786 358787 14789
rect 111425 14784 358787 14786
rect 111425 14728 111430 14784
rect 111486 14728 358726 14784
rect 358782 14728 358787 14784
rect 111425 14726 358787 14728
rect 96337 14723 96403 14726
rect 111425 14723 111491 14726
rect 358721 14723 358787 14726
rect 19926 14588 19932 14652
rect 19996 14650 20002 14652
rect 92565 14650 92631 14653
rect 19996 14648 92631 14650
rect 19996 14592 92570 14648
rect 92626 14592 92631 14648
rect 19996 14590 92631 14592
rect 19996 14588 20002 14590
rect 92565 14587 92631 14590
rect 97165 14650 97231 14653
rect 367645 14650 367711 14653
rect 97165 14648 367711 14650
rect 97165 14592 97170 14648
rect 97226 14592 367650 14648
rect 367706 14592 367711 14648
rect 97165 14590 367711 14592
rect 97165 14587 97231 14590
rect 367645 14587 367711 14590
rect 15009 14514 15075 14517
rect 96521 14514 96587 14517
rect 15009 14512 96587 14514
rect 15009 14456 15014 14512
rect 15070 14456 96526 14512
rect 96582 14456 96587 14512
rect 15009 14454 96587 14456
rect 15009 14451 15075 14454
rect 96521 14451 96587 14454
rect 97073 14514 97139 14517
rect 104801 14514 104867 14517
rect 97073 14512 104867 14514
rect 97073 14456 97078 14512
rect 97134 14456 104806 14512
rect 104862 14456 104867 14512
rect 97073 14454 104867 14456
rect 97073 14451 97139 14454
rect 104801 14451 104867 14454
rect 113817 14514 113883 14517
rect 430573 14514 430639 14517
rect 113817 14512 430639 14514
rect 113817 14456 113822 14512
rect 113878 14456 430578 14512
rect 430634 14456 430639 14512
rect 113817 14454 430639 14456
rect 113817 14451 113883 14454
rect 430573 14451 430639 14454
rect 116117 14106 116183 14109
rect 118785 14106 118851 14109
rect 116117 14104 118851 14106
rect 116117 14048 116122 14104
rect 116178 14048 118790 14104
rect 118846 14048 118851 14104
rect 116117 14046 118851 14048
rect 116117 14043 116183 14046
rect 118785 14043 118851 14046
rect 124213 13970 124279 13973
rect 124213 13968 129842 13970
rect 124213 13912 124218 13968
rect 124274 13912 129842 13968
rect 124213 13910 129842 13912
rect 124213 13907 124279 13910
rect 94405 13834 94471 13837
rect 96889 13834 96955 13837
rect 94405 13832 96955 13834
rect 94405 13776 94410 13832
rect 94466 13776 96894 13832
rect 96950 13776 96955 13832
rect 94405 13774 96955 13776
rect 94405 13771 94471 13774
rect 96889 13771 96955 13774
rect 117037 13834 117103 13837
rect 123661 13834 123727 13837
rect 124213 13834 124279 13837
rect 117037 13832 118618 13834
rect 117037 13776 117042 13832
rect 117098 13776 118618 13832
rect 117037 13774 118618 13776
rect 117037 13771 117103 13774
rect 59169 13698 59235 13701
rect 96337 13698 96403 13701
rect 59169 13696 96403 13698
rect 59169 13640 59174 13696
rect 59230 13640 96342 13696
rect 96398 13640 96403 13696
rect 59169 13638 96403 13640
rect 59169 13635 59235 13638
rect 96337 13635 96403 13638
rect 96521 13698 96587 13701
rect 105813 13698 105879 13701
rect 96521 13696 105879 13698
rect 96521 13640 96526 13696
rect 96582 13640 105818 13696
rect 105874 13640 105879 13696
rect 96521 13638 105879 13640
rect 96521 13635 96587 13638
rect 105813 13635 105879 13638
rect 114369 13698 114435 13701
rect 118325 13698 118391 13701
rect 114369 13696 118391 13698
rect 114369 13640 114374 13696
rect 114430 13640 118330 13696
rect 118386 13640 118391 13696
rect 114369 13638 118391 13640
rect 114369 13635 114435 13638
rect 118325 13635 118391 13638
rect 95785 13562 95851 13565
rect 97809 13562 97875 13565
rect 95785 13560 97875 13562
rect 95785 13504 95790 13560
rect 95846 13504 97814 13560
rect 97870 13504 97875 13560
rect 95785 13502 97875 13504
rect 95785 13499 95851 13502
rect 97809 13499 97875 13502
rect 114461 13562 114527 13565
rect 114737 13562 114803 13565
rect 114461 13560 114803 13562
rect 114461 13504 114466 13560
rect 114522 13504 114742 13560
rect 114798 13504 114803 13560
rect 114461 13502 114803 13504
rect 114461 13499 114527 13502
rect 114737 13499 114803 13502
rect 117221 13562 117287 13565
rect 118233 13562 118299 13565
rect 117221 13560 118299 13562
rect 117221 13504 117226 13560
rect 117282 13504 118238 13560
rect 118294 13504 118299 13560
rect 117221 13502 118299 13504
rect 118558 13562 118618 13774
rect 123661 13832 124279 13834
rect 123661 13776 123666 13832
rect 123722 13776 124218 13832
rect 124274 13776 124279 13832
rect 123661 13774 124279 13776
rect 123661 13771 123727 13774
rect 124213 13771 124279 13774
rect 125869 13834 125935 13837
rect 128997 13834 129063 13837
rect 125869 13832 129063 13834
rect 125869 13776 125874 13832
rect 125930 13776 129002 13832
rect 129058 13776 129063 13832
rect 125869 13774 129063 13776
rect 125869 13771 125935 13774
rect 128997 13771 129063 13774
rect 129782 13698 129842 13910
rect 132585 13698 132651 13701
rect 129782 13696 132651 13698
rect 129782 13640 132590 13696
rect 132646 13640 132651 13696
rect 129782 13638 132651 13640
rect 132585 13635 132651 13638
rect 137277 13698 137343 13701
rect 155493 13698 155559 13701
rect 137277 13696 155559 13698
rect 137277 13640 137282 13696
rect 137338 13640 155498 13696
rect 155554 13640 155559 13696
rect 137277 13638 155559 13640
rect 137277 13635 137343 13638
rect 155493 13635 155559 13638
rect 150525 13562 150591 13565
rect 118558 13560 150591 13562
rect 118558 13504 150530 13560
rect 150586 13504 150591 13560
rect 118558 13502 150591 13504
rect 117221 13499 117287 13502
rect 118233 13499 118299 13502
rect 150525 13499 150591 13502
rect 107561 13426 107627 13429
rect 122833 13426 122899 13429
rect 107561 13424 122899 13426
rect 107561 13368 107566 13424
rect 107622 13368 122838 13424
rect 122894 13368 122899 13424
rect 107561 13366 122899 13368
rect 107561 13363 107627 13366
rect 122833 13363 122899 13366
rect 125317 13426 125383 13429
rect 154297 13426 154363 13429
rect 125317 13424 154363 13426
rect 125317 13368 125322 13424
rect 125378 13368 154302 13424
rect 154358 13368 154363 13424
rect 125317 13366 154363 13368
rect 125317 13363 125383 13366
rect 154297 13363 154363 13366
rect 98177 13290 98243 13293
rect 371233 13290 371299 13293
rect 98177 13288 371299 13290
rect 98177 13232 98182 13288
rect 98238 13232 371238 13288
rect 371294 13232 371299 13288
rect 98177 13230 371299 13232
rect 98177 13227 98243 13230
rect 371233 13227 371299 13230
rect 22093 13154 22159 13157
rect 107561 13154 107627 13157
rect 420913 13154 420979 13157
rect 22093 13152 107627 13154
rect 22093 13096 22098 13152
rect 22154 13096 107566 13152
rect 107622 13096 107627 13152
rect 22093 13094 107627 13096
rect 22093 13091 22159 13094
rect 107561 13091 107627 13094
rect 107702 13152 420979 13154
rect 107702 13096 420918 13152
rect 420974 13096 420979 13152
rect 107702 13094 420979 13096
rect 12341 13018 12407 13021
rect 96521 13018 96587 13021
rect 12341 13016 96587 13018
rect 12341 12960 12346 13016
rect 12402 12960 96526 13016
rect 96582 12960 96587 13016
rect 12341 12958 96587 12960
rect 12341 12955 12407 12958
rect 96521 12955 96587 12958
rect 105445 13018 105511 13021
rect 107702 13018 107762 13094
rect 420913 13091 420979 13094
rect 105445 13016 107762 13018
rect 105445 12960 105450 13016
rect 105506 12960 107762 13016
rect 105445 12958 107762 12960
rect 117497 13018 117563 13021
rect 482369 13018 482435 13021
rect 117497 13016 482435 13018
rect 117497 12960 117502 13016
rect 117558 12960 482374 13016
rect 482430 12960 482435 13016
rect 117497 12958 482435 12960
rect 105445 12955 105511 12958
rect 117497 12955 117563 12958
rect 482369 12955 482435 12958
rect 104157 12882 104223 12885
rect 114185 12882 114251 12885
rect 104157 12880 114251 12882
rect 104157 12824 104162 12880
rect 104218 12824 114190 12880
rect 114246 12824 114251 12880
rect 104157 12822 114251 12824
rect 104157 12819 104223 12822
rect 114185 12819 114251 12822
rect 121361 12746 121427 12749
rect 157333 12746 157399 12749
rect 121361 12744 157399 12746
rect 121361 12688 121366 12744
rect 121422 12688 157338 12744
rect 157394 12688 157399 12744
rect 121361 12686 157399 12688
rect 121361 12683 121427 12686
rect 157333 12683 157399 12686
rect 95141 12474 95207 12477
rect 115933 12474 115999 12477
rect 118601 12474 118667 12477
rect 95141 12472 98010 12474
rect 95141 12416 95146 12472
rect 95202 12416 98010 12472
rect 95141 12414 98010 12416
rect 95141 12411 95207 12414
rect 19149 12338 19215 12341
rect 94957 12338 95023 12341
rect 19149 12336 95023 12338
rect 19149 12280 19154 12336
rect 19210 12280 94962 12336
rect 95018 12280 95023 12336
rect 19149 12278 95023 12280
rect 97950 12338 98010 12414
rect 115933 12472 118667 12474
rect 115933 12416 115938 12472
rect 115994 12416 118606 12472
rect 118662 12416 118667 12472
rect 115933 12414 118667 12416
rect 115933 12411 115999 12414
rect 118601 12411 118667 12414
rect 107745 12338 107811 12341
rect 97950 12336 107811 12338
rect 97950 12280 107750 12336
rect 107806 12280 107811 12336
rect 97950 12278 107811 12280
rect 19149 12275 19215 12278
rect 94957 12275 95023 12278
rect 107745 12275 107811 12278
rect 111149 12338 111215 12341
rect 114461 12338 114527 12341
rect 111149 12336 114527 12338
rect 111149 12280 111154 12336
rect 111210 12280 114466 12336
rect 114522 12280 114527 12336
rect 111149 12278 114527 12280
rect 111149 12275 111215 12278
rect 114461 12275 114527 12278
rect 96521 12202 96587 12205
rect 100845 12202 100911 12205
rect 96521 12200 100911 12202
rect 96521 12144 96526 12200
rect 96582 12144 100850 12200
rect 100906 12144 100911 12200
rect 96521 12142 100911 12144
rect 96521 12139 96587 12142
rect 100845 12139 100911 12142
rect 119981 12202 120047 12205
rect 150893 12202 150959 12205
rect 119981 12200 150959 12202
rect 119981 12144 119986 12200
rect 120042 12144 150898 12200
rect 150954 12144 150959 12200
rect 119981 12142 150959 12144
rect 119981 12139 120047 12142
rect 150893 12139 150959 12142
rect 107469 12066 107535 12069
rect 126237 12066 126303 12069
rect 155953 12066 156019 12069
rect 107469 12064 113190 12066
rect 107469 12008 107474 12064
rect 107530 12008 113190 12064
rect 107469 12006 113190 12008
rect 107469 12003 107535 12006
rect 84377 11930 84443 11933
rect 95233 11930 95299 11933
rect 84377 11928 95299 11930
rect 84377 11872 84382 11928
rect 84438 11872 95238 11928
rect 95294 11872 95299 11928
rect 84377 11870 95299 11872
rect 84377 11867 84443 11870
rect 95233 11867 95299 11870
rect 101489 11930 101555 11933
rect 107561 11930 107627 11933
rect 101489 11928 107627 11930
rect 101489 11872 101494 11928
rect 101550 11872 107566 11928
rect 107622 11872 107627 11928
rect 101489 11870 107627 11872
rect 113130 11930 113190 12006
rect 126237 12064 156019 12066
rect 126237 12008 126242 12064
rect 126298 12008 155958 12064
rect 156014 12008 156019 12064
rect 126237 12006 156019 12008
rect 126237 12003 126303 12006
rect 155953 12003 156019 12006
rect 377949 11930 378015 11933
rect 113130 11928 378015 11930
rect 113130 11872 377954 11928
rect 378010 11872 378015 11928
rect 113130 11870 378015 11872
rect 101489 11867 101555 11870
rect 107561 11867 107627 11870
rect 377949 11867 378015 11870
rect 82445 11794 82511 11797
rect 102409 11794 102475 11797
rect 82445 11792 102475 11794
rect 82445 11736 82450 11792
rect 82506 11736 102414 11792
rect 102470 11736 102475 11792
rect 82445 11734 102475 11736
rect 82445 11731 82511 11734
rect 102409 11731 102475 11734
rect 108573 11794 108639 11797
rect 404261 11794 404327 11797
rect 108573 11792 404327 11794
rect 108573 11736 108578 11792
rect 108634 11736 404266 11792
rect 404322 11736 404327 11792
rect 108573 11734 404327 11736
rect 108573 11731 108639 11734
rect 404261 11731 404327 11734
rect 35985 11658 36051 11661
rect 83181 11658 83247 11661
rect 35985 11656 83247 11658
rect 35985 11600 35990 11656
rect 36046 11600 83186 11656
rect 83242 11600 83247 11656
rect 35985 11598 83247 11600
rect 35985 11595 36051 11598
rect 83181 11595 83247 11598
rect 92565 11658 92631 11661
rect 106089 11658 106155 11661
rect 92565 11656 106155 11658
rect 92565 11600 92570 11656
rect 92626 11600 106094 11656
rect 106150 11600 106155 11656
rect 92565 11598 106155 11600
rect 92565 11595 92631 11598
rect 106089 11595 106155 11598
rect 110413 11658 110479 11661
rect 453205 11658 453271 11661
rect 110413 11656 453271 11658
rect 110413 11600 110418 11656
rect 110474 11600 453210 11656
rect 453266 11600 453271 11656
rect 110413 11598 453271 11600
rect 110413 11595 110479 11598
rect 453205 11595 453271 11598
rect 114093 11522 114159 11525
rect 126881 11522 126947 11525
rect 154113 11522 154179 11525
rect 114093 11520 122850 11522
rect 114093 11464 114098 11520
rect 114154 11464 122850 11520
rect 114093 11462 122850 11464
rect 114093 11459 114159 11462
rect 112621 11386 112687 11389
rect 115749 11386 115815 11389
rect 112621 11384 115815 11386
rect 112621 11328 112626 11384
rect 112682 11328 115754 11384
rect 115810 11328 115815 11384
rect 112621 11326 115815 11328
rect 122790 11386 122850 11462
rect 126881 11520 154179 11522
rect 126881 11464 126886 11520
rect 126942 11464 154118 11520
rect 154174 11464 154179 11520
rect 126881 11462 154179 11464
rect 126881 11459 126947 11462
rect 154113 11459 154179 11462
rect 149053 11386 149119 11389
rect 122790 11384 149119 11386
rect 122790 11328 149058 11384
rect 149114 11328 149119 11384
rect 122790 11326 149119 11328
rect 112621 11323 112687 11326
rect 115749 11323 115815 11326
rect 149053 11323 149119 11326
rect 105629 11250 105695 11253
rect 110505 11250 110571 11253
rect 105629 11248 110571 11250
rect 105629 11192 105634 11248
rect 105690 11192 110510 11248
rect 110566 11192 110571 11248
rect 105629 11190 110571 11192
rect 105629 11187 105695 11190
rect 110505 11187 110571 11190
rect 111609 11114 111675 11117
rect 124121 11114 124187 11117
rect 111609 11112 111810 11114
rect 111609 11056 111614 11112
rect 111670 11056 111810 11112
rect 111609 11054 111810 11056
rect 111609 11051 111675 11054
rect 21357 10978 21423 10981
rect 98085 10978 98151 10981
rect 21357 10976 98151 10978
rect 21357 10920 21362 10976
rect 21418 10920 98090 10976
rect 98146 10920 98151 10976
rect 21357 10918 98151 10920
rect 111750 10978 111810 11054
rect 124121 11112 127082 11114
rect 124121 11056 124126 11112
rect 124182 11056 127082 11112
rect 124121 11054 127082 11056
rect 124121 11051 124187 11054
rect 115749 10978 115815 10981
rect 111750 10976 115815 10978
rect 111750 10920 115754 10976
rect 115810 10920 115815 10976
rect 111750 10918 115815 10920
rect 21357 10915 21423 10918
rect 98085 10915 98151 10918
rect 115749 10915 115815 10918
rect 119245 10978 119311 10981
rect 126881 10978 126947 10981
rect 119245 10976 126947 10978
rect 119245 10920 119250 10976
rect 119306 10920 126886 10976
rect 126942 10920 126947 10976
rect 119245 10918 126947 10920
rect 127022 10978 127082 11054
rect 133229 10978 133295 10981
rect 156689 10978 156755 10981
rect 127022 10976 133295 10978
rect 127022 10920 133234 10976
rect 133290 10920 133295 10976
rect 127022 10918 133295 10920
rect 119245 10915 119311 10918
rect 126881 10915 126947 10918
rect 133229 10915 133295 10918
rect 142110 10976 156755 10978
rect 142110 10920 156694 10976
rect 156750 10920 156755 10976
rect 142110 10918 156755 10920
rect 77201 10842 77267 10845
rect 95785 10842 95851 10845
rect 77201 10840 95851 10842
rect 77201 10784 77206 10840
rect 77262 10784 95790 10840
rect 95846 10784 95851 10840
rect 77201 10782 95851 10784
rect 77201 10779 77267 10782
rect 95785 10779 95851 10782
rect 107377 10842 107443 10845
rect 117589 10842 117655 10845
rect 107377 10840 117655 10842
rect 107377 10784 107382 10840
rect 107438 10784 117594 10840
rect 117650 10784 117655 10840
rect 107377 10782 117655 10784
rect 107377 10779 107443 10782
rect 117589 10779 117655 10782
rect 128905 10842 128971 10845
rect 142110 10842 142170 10918
rect 156689 10915 156755 10918
rect 128905 10840 142170 10842
rect 128905 10784 128910 10840
rect 128966 10784 142170 10840
rect 128905 10782 142170 10784
rect 128905 10779 128971 10782
rect 79225 10706 79291 10709
rect 104525 10706 104591 10709
rect 79225 10704 104591 10706
rect 79225 10648 79230 10704
rect 79286 10648 104530 10704
rect 104586 10648 104591 10704
rect 79225 10646 104591 10648
rect 79225 10643 79291 10646
rect 104525 10643 104591 10646
rect 100293 10570 100359 10573
rect 377397 10570 377463 10573
rect 100293 10568 377463 10570
rect 100293 10512 100298 10568
rect 100354 10512 377402 10568
rect 377458 10512 377463 10568
rect 100293 10510 377463 10512
rect 100293 10507 100359 10510
rect 377397 10507 377463 10510
rect 102501 10434 102567 10437
rect 385309 10434 385375 10437
rect 102501 10432 385375 10434
rect 102501 10376 102506 10432
rect 102562 10376 385314 10432
rect 385370 10376 385375 10432
rect 102501 10374 385375 10376
rect 102501 10371 102567 10374
rect 385309 10371 385375 10374
rect 23105 10298 23171 10301
rect 88425 10298 88491 10301
rect 23105 10296 88491 10298
rect 23105 10240 23110 10296
rect 23166 10240 88430 10296
rect 88486 10240 88491 10296
rect 23105 10238 88491 10240
rect 23105 10235 23171 10238
rect 88425 10235 88491 10238
rect 95233 10298 95299 10301
rect 104801 10298 104867 10301
rect 95233 10296 104867 10298
rect 95233 10240 95238 10296
rect 95294 10240 104806 10296
rect 104862 10240 104867 10296
rect 95233 10238 104867 10240
rect 95233 10235 95299 10238
rect 104801 10235 104867 10238
rect 109033 10298 109099 10301
rect 442625 10298 442691 10301
rect 109033 10296 442691 10298
rect 109033 10240 109038 10296
rect 109094 10240 442630 10296
rect 442686 10240 442691 10296
rect 109033 10238 442691 10240
rect 109033 10235 109099 10238
rect 442625 10235 442691 10238
rect 106089 9754 106155 9757
rect 119889 9754 119955 9757
rect 106089 9752 106290 9754
rect 106089 9696 106094 9752
rect 106150 9696 106290 9752
rect 106089 9694 106290 9696
rect 106089 9691 106155 9694
rect 10961 9618 11027 9621
rect 106230 9618 106290 9694
rect 119889 9752 132510 9754
rect 119889 9696 119894 9752
rect 119950 9696 132510 9752
rect 119889 9694 132510 9696
rect 119889 9691 119955 9694
rect 110597 9618 110663 9621
rect 10961 9616 103530 9618
rect 10961 9560 10966 9616
rect 11022 9560 103530 9616
rect 10961 9558 103530 9560
rect 106230 9616 110663 9618
rect 106230 9560 110602 9616
rect 110658 9560 110663 9616
rect 106230 9558 110663 9560
rect 10961 9555 11027 9558
rect 23749 9482 23815 9485
rect 98729 9482 98795 9485
rect 23749 9480 98795 9482
rect 23749 9424 23754 9480
rect 23810 9424 98734 9480
rect 98790 9424 98795 9480
rect 23749 9422 98795 9424
rect 103470 9482 103530 9558
rect 110597 9555 110663 9558
rect 113357 9618 113423 9621
rect 120073 9618 120139 9621
rect 113357 9616 120139 9618
rect 113357 9560 113362 9616
rect 113418 9560 120078 9616
rect 120134 9560 120139 9616
rect 113357 9558 120139 9560
rect 132450 9618 132510 9694
rect 152549 9618 152615 9621
rect 132450 9616 152615 9618
rect 132450 9560 152554 9616
rect 152610 9560 152615 9616
rect 132450 9558 152615 9560
rect 113357 9555 113423 9558
rect 120073 9555 120139 9558
rect 152549 9555 152615 9558
rect 111977 9482 112043 9485
rect 103470 9480 112043 9482
rect 103470 9424 111982 9480
rect 112038 9424 112043 9480
rect 103470 9422 112043 9424
rect 23749 9419 23815 9422
rect 98729 9419 98795 9422
rect 111977 9419 112043 9422
rect 121269 9482 121335 9485
rect 151169 9482 151235 9485
rect 121269 9480 151235 9482
rect 121269 9424 121274 9480
rect 121330 9424 151174 9480
rect 151230 9424 151235 9480
rect 121269 9422 151235 9424
rect 121269 9419 121335 9422
rect 151169 9419 151235 9422
rect 91185 9346 91251 9349
rect 114369 9346 114435 9349
rect 91185 9344 114435 9346
rect 91185 9288 91190 9344
rect 91246 9288 114374 9344
rect 114430 9288 114435 9344
rect 91185 9286 114435 9288
rect 91185 9283 91251 9286
rect 114369 9283 114435 9286
rect 117129 9346 117195 9349
rect 403709 9346 403775 9349
rect 117129 9344 403775 9346
rect 117129 9288 117134 9344
rect 117190 9288 403714 9344
rect 403770 9288 403775 9344
rect 117129 9286 403775 9288
rect 117129 9283 117195 9286
rect 403709 9283 403775 9286
rect 104341 9210 104407 9213
rect 414289 9210 414355 9213
rect 104341 9208 414355 9210
rect 104341 9152 104346 9208
rect 104402 9152 414294 9208
rect 414350 9152 414355 9208
rect 104341 9150 414355 9152
rect 104341 9147 104407 9150
rect 414289 9147 414355 9150
rect 113173 9074 113239 9077
rect 462313 9074 462379 9077
rect 113173 9072 462379 9074
rect 113173 9016 113178 9072
rect 113234 9016 462318 9072
rect 462374 9016 462379 9072
rect 113173 9014 462379 9016
rect 113173 9011 113239 9014
rect 462313 9011 462379 9014
rect 88425 8938 88491 8941
rect 101397 8938 101463 8941
rect 88425 8936 101463 8938
rect 88425 8880 88430 8936
rect 88486 8880 101402 8936
rect 101458 8880 101463 8936
rect 88425 8878 101463 8880
rect 88425 8875 88491 8878
rect 101397 8875 101463 8878
rect 124213 8938 124279 8941
rect 538397 8938 538463 8941
rect 124213 8936 538463 8938
rect 124213 8880 124218 8936
rect 124274 8880 538402 8936
rect 538458 8880 538463 8936
rect 124213 8878 538463 8880
rect 124213 8875 124279 8878
rect 538397 8875 538463 8878
rect 140773 8802 140839 8805
rect 154113 8802 154179 8805
rect 140773 8800 154179 8802
rect 140773 8744 140778 8800
rect 140834 8744 154118 8800
rect 154174 8744 154179 8800
rect 140773 8742 154179 8744
rect 140773 8739 140839 8742
rect 154113 8739 154179 8742
rect 110505 8394 110571 8397
rect 113173 8394 113239 8397
rect 110505 8392 113239 8394
rect 110505 8336 110510 8392
rect 110566 8336 113178 8392
rect 113234 8336 113239 8392
rect 110505 8334 113239 8336
rect 110505 8331 110571 8334
rect 113173 8331 113239 8334
rect 63585 8258 63651 8261
rect 104249 8258 104315 8261
rect 63585 8256 104315 8258
rect 63585 8200 63590 8256
rect 63646 8200 104254 8256
rect 104310 8200 104315 8256
rect 63585 8198 104315 8200
rect 63585 8195 63651 8198
rect 104249 8195 104315 8198
rect 114645 8258 114711 8261
rect 353017 8258 353083 8261
rect 114645 8256 353083 8258
rect 114645 8200 114650 8256
rect 114706 8200 353022 8256
rect 353078 8200 353083 8256
rect 114645 8198 353083 8200
rect 114645 8195 114711 8198
rect 353017 8195 353083 8198
rect 71773 8122 71839 8125
rect 97993 8122 98059 8125
rect 71773 8120 98059 8122
rect 71773 8064 71778 8120
rect 71834 8064 97998 8120
rect 98054 8064 98059 8120
rect 71773 8062 98059 8064
rect 71773 8059 71839 8062
rect 97993 8059 98059 8062
rect 105997 8122 106063 8125
rect 424961 8122 425027 8125
rect 105997 8120 425027 8122
rect 105997 8064 106002 8120
rect 106058 8064 424966 8120
rect 425022 8064 425027 8120
rect 105997 8062 425027 8064
rect 105997 8059 106063 8062
rect 424961 8059 425027 8062
rect 86953 7986 87019 7989
rect 102133 7986 102199 7989
rect 86953 7984 102199 7986
rect 86953 7928 86958 7984
rect 87014 7928 102138 7984
rect 102194 7928 102199 7984
rect 86953 7926 102199 7928
rect 86953 7923 87019 7926
rect 102133 7923 102199 7926
rect 106549 7986 106615 7989
rect 428457 7986 428523 7989
rect 106549 7984 428523 7986
rect 106549 7928 106554 7984
rect 106610 7928 428462 7984
rect 428518 7928 428523 7984
rect 106549 7926 428523 7928
rect 106549 7923 106615 7926
rect 428457 7923 428523 7926
rect 115565 7850 115631 7853
rect 486417 7850 486483 7853
rect 115565 7848 486483 7850
rect 115565 7792 115570 7848
rect 115626 7792 486422 7848
rect 486478 7792 486483 7848
rect 115565 7790 486483 7792
rect 115565 7787 115631 7790
rect 486417 7787 486483 7790
rect 104893 7714 104959 7717
rect 114829 7714 114895 7717
rect 104893 7712 114895 7714
rect 104893 7656 104898 7712
rect 104954 7656 114834 7712
rect 114890 7656 114895 7712
rect 104893 7654 114895 7656
rect 104893 7651 104959 7654
rect 114829 7651 114895 7654
rect 120533 7714 120599 7717
rect 518341 7714 518407 7717
rect 120533 7712 518407 7714
rect 120533 7656 120538 7712
rect 120594 7656 518346 7712
rect 518402 7656 518407 7712
rect 120533 7654 518407 7656
rect 120533 7651 120599 7654
rect 518341 7651 518407 7654
rect 97993 7578 98059 7581
rect 115841 7578 115907 7581
rect 97993 7576 115907 7578
rect 97993 7520 97998 7576
rect 98054 7520 115846 7576
rect 115902 7520 115907 7576
rect 97993 7518 115907 7520
rect 97993 7515 98059 7518
rect 115841 7515 115907 7518
rect 127709 7578 127775 7581
rect 562317 7578 562383 7581
rect 127709 7576 562383 7578
rect 127709 7520 127714 7576
rect 127770 7520 562322 7576
rect 562378 7520 562383 7576
rect 127709 7518 562383 7520
rect 127709 7515 127775 7518
rect 562317 7515 562383 7518
rect 108021 7306 108087 7309
rect 114461 7306 114527 7309
rect 108021 7304 114527 7306
rect 108021 7248 108026 7304
rect 108082 7248 114466 7304
rect 114522 7248 114527 7304
rect 108021 7246 114527 7248
rect 108021 7243 108087 7246
rect 114461 7243 114527 7246
rect 102133 7034 102199 7037
rect 107561 7034 107627 7037
rect 102133 7032 107627 7034
rect 102133 6976 102138 7032
rect 102194 6976 107566 7032
rect 107622 6976 107627 7032
rect 102133 6974 107627 6976
rect 102133 6971 102199 6974
rect 107561 6971 107627 6974
rect 35893 6898 35959 6901
rect 97993 6898 98059 6901
rect 35893 6896 98059 6898
rect 35893 6840 35898 6896
rect 35954 6840 97998 6896
rect 98054 6840 98059 6896
rect 35893 6838 98059 6840
rect 35893 6835 35959 6838
rect 97993 6835 98059 6838
rect 104525 6898 104591 6901
rect 108389 6898 108455 6901
rect 104525 6896 108455 6898
rect 104525 6840 104530 6896
rect 104586 6840 108394 6896
rect 108450 6840 108455 6896
rect 104525 6838 108455 6840
rect 104525 6835 104591 6838
rect 108389 6835 108455 6838
rect 115289 6898 115355 6901
rect 118693 6898 118759 6901
rect 115289 6896 118759 6898
rect 115289 6840 115294 6896
rect 115350 6840 118698 6896
rect 118754 6840 118759 6896
rect 115289 6838 118759 6840
rect 115289 6835 115355 6838
rect 118693 6835 118759 6838
rect 96245 6762 96311 6765
rect 358813 6762 358879 6765
rect 96245 6760 358879 6762
rect 96245 6704 96250 6760
rect 96306 6704 358818 6760
rect 358874 6704 358879 6760
rect 96245 6702 358879 6704
rect 96245 6699 96311 6702
rect 358813 6699 358879 6702
rect 82077 6626 82143 6629
rect 96797 6626 96863 6629
rect 82077 6624 96863 6626
rect -960 6490 480 6580
rect 82077 6568 82082 6624
rect 82138 6568 96802 6624
rect 96858 6568 96863 6624
rect 82077 6566 96863 6568
rect 82077 6563 82143 6566
rect 96797 6563 96863 6566
rect 98453 6626 98519 6629
rect 372613 6626 372679 6629
rect 98453 6624 372679 6626
rect 98453 6568 98458 6624
rect 98514 6568 372618 6624
rect 372674 6568 372679 6624
rect 98453 6566 372679 6568
rect 98453 6563 98519 6566
rect 372613 6563 372679 6566
rect 578877 6626 578943 6629
rect 583520 6626 584960 6716
rect 578877 6624 584960 6626
rect 578877 6568 578882 6624
rect 578938 6568 584960 6624
rect 578877 6566 584960 6568
rect 578877 6563 578943 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 98821 6490 98887 6493
rect 378869 6490 378935 6493
rect 98821 6488 378935 6490
rect 98821 6432 98826 6488
rect 98882 6432 378874 6488
rect 378930 6432 378935 6488
rect 583520 6476 584960 6566
rect 98821 6430 378935 6432
rect 98821 6427 98887 6430
rect 378869 6427 378935 6430
rect 103237 6354 103303 6357
rect 407205 6354 407271 6357
rect 103237 6352 407271 6354
rect 103237 6296 103242 6352
rect 103298 6296 407210 6352
rect 407266 6296 407271 6352
rect 103237 6294 407271 6296
rect 103237 6291 103303 6294
rect 407205 6291 407271 6294
rect 33869 6218 33935 6221
rect 95233 6218 95299 6221
rect 33869 6216 95299 6218
rect 33869 6160 33874 6216
rect 33930 6160 95238 6216
rect 95294 6160 95299 6216
rect 33869 6158 95299 6160
rect 33869 6155 33935 6158
rect 95233 6155 95299 6158
rect 107653 6218 107719 6221
rect 435541 6218 435607 6221
rect 107653 6216 435607 6218
rect 107653 6160 107658 6216
rect 107714 6160 435546 6216
rect 435602 6160 435607 6216
rect 107653 6158 435607 6160
rect 107653 6155 107719 6158
rect 435541 6155 435607 6158
rect 70669 6082 70735 6085
rect 102133 6082 102199 6085
rect 70669 6080 102199 6082
rect 70669 6024 70674 6080
rect 70730 6024 102138 6080
rect 102194 6024 102199 6080
rect 70669 6022 102199 6024
rect 70669 6019 70735 6022
rect 102133 6019 102199 6022
rect 110597 6082 110663 6085
rect 114461 6082 114527 6085
rect 110597 6080 114527 6082
rect 110597 6024 110602 6080
rect 110658 6024 114466 6080
rect 114522 6024 114527 6080
rect 110597 6022 114527 6024
rect 110597 6019 110663 6022
rect 114461 6019 114527 6022
rect 140681 6082 140747 6085
rect 147029 6082 147095 6085
rect 140681 6080 147095 6082
rect 140681 6024 140686 6080
rect 140742 6024 147034 6080
rect 147090 6024 147095 6080
rect 140681 6022 147095 6024
rect 140681 6019 140747 6022
rect 147029 6019 147095 6022
rect 113173 5946 113239 5949
rect 120809 5946 120875 5949
rect 113173 5944 120875 5946
rect 113173 5888 113178 5944
rect 113234 5888 120814 5944
rect 120870 5888 120875 5944
rect 113173 5886 120875 5888
rect 113173 5883 113239 5886
rect 120809 5883 120875 5886
rect 130653 5674 130719 5677
rect 143533 5674 143599 5677
rect 130653 5672 143599 5674
rect 130653 5616 130658 5672
rect 130714 5616 143538 5672
rect 143594 5616 143599 5672
rect 130653 5614 143599 5616
rect 130653 5611 130719 5614
rect 143533 5611 143599 5614
rect 97625 5538 97691 5541
rect 329189 5538 329255 5541
rect 97625 5536 329255 5538
rect 97625 5480 97630 5536
rect 97686 5480 329194 5536
rect 329250 5480 329255 5536
rect 97625 5478 329255 5480
rect 97625 5475 97691 5478
rect 329189 5475 329255 5478
rect 95049 5402 95115 5405
rect 340965 5402 341031 5405
rect 95049 5400 341031 5402
rect 95049 5344 95054 5400
rect 95110 5344 340970 5400
rect 341026 5344 341031 5400
rect 95049 5342 341031 5344
rect 95049 5339 95115 5342
rect 340965 5339 341031 5342
rect 100477 5266 100543 5269
rect 389449 5266 389515 5269
rect 100477 5264 389515 5266
rect 100477 5208 100482 5264
rect 100538 5208 389454 5264
rect 389510 5208 389515 5264
rect 100477 5206 389515 5208
rect 100477 5203 100543 5206
rect 389449 5203 389515 5206
rect 81341 5130 81407 5133
rect 104157 5130 104223 5133
rect 81341 5128 104223 5130
rect 81341 5072 81346 5128
rect 81402 5072 104162 5128
rect 104218 5072 104223 5128
rect 81341 5070 104223 5072
rect 81341 5067 81407 5070
rect 104157 5067 104223 5070
rect 108205 5130 108271 5133
rect 439129 5130 439195 5133
rect 108205 5128 439195 5130
rect 108205 5072 108210 5128
rect 108266 5072 439134 5128
rect 439190 5072 439195 5128
rect 108205 5070 439195 5072
rect 108205 5067 108271 5070
rect 439129 5067 439195 5070
rect 121637 4994 121703 4997
rect 525425 4994 525491 4997
rect 121637 4992 525491 4994
rect 121637 4936 121642 4992
rect 121698 4936 525430 4992
rect 525486 4936 525491 4992
rect 121637 4934 525491 4936
rect 121637 4931 121703 4934
rect 525425 4931 525491 4934
rect 71037 4858 71103 4861
rect 104433 4858 104499 4861
rect 71037 4856 104499 4858
rect 71037 4800 71042 4856
rect 71098 4800 104438 4856
rect 104494 4800 104499 4856
rect 71037 4798 104499 4800
rect 71037 4795 71103 4798
rect 104433 4795 104499 4798
rect 129917 4858 129983 4861
rect 578601 4858 578667 4861
rect 129917 4856 578667 4858
rect 129917 4800 129922 4856
rect 129978 4800 578606 4856
rect 578662 4800 578667 4856
rect 129917 4798 578667 4800
rect 129917 4795 129983 4798
rect 578601 4795 578667 4798
rect 128997 4722 129063 4725
rect 146937 4722 147003 4725
rect 128997 4720 147003 4722
rect 128997 4664 129002 4720
rect 129058 4664 146942 4720
rect 146998 4664 147003 4720
rect 128997 4662 147003 4664
rect 128997 4659 129063 4662
rect 146937 4659 147003 4662
rect 103513 4314 103579 4317
rect 108021 4314 108087 4317
rect 103513 4312 108087 4314
rect 103513 4256 103518 4312
rect 103574 4256 108026 4312
rect 108082 4256 108087 4312
rect 103513 4254 108087 4256
rect 103513 4251 103579 4254
rect 108021 4251 108087 4254
rect 101765 4178 101831 4181
rect 101765 4176 103714 4178
rect 101765 4120 101770 4176
rect 101826 4120 103714 4176
rect 101765 4118 103714 4120
rect 101765 4115 101831 4118
rect 88333 4042 88399 4045
rect 103513 4042 103579 4045
rect 88333 4040 103579 4042
rect 88333 3984 88338 4040
rect 88394 3984 103518 4040
rect 103574 3984 103579 4040
rect 88333 3982 103579 3984
rect 103654 4042 103714 4118
rect 150433 4042 150499 4045
rect 103654 4040 150499 4042
rect 103654 3984 150438 4040
rect 150494 3984 150499 4040
rect 103654 3982 150499 3984
rect 88333 3979 88399 3982
rect 103513 3979 103579 3982
rect 150433 3979 150499 3982
rect 114093 3906 114159 3909
rect 122373 3906 122439 3909
rect 114093 3904 122439 3906
rect 114093 3848 114098 3904
rect 114154 3848 122378 3904
rect 122434 3848 122439 3904
rect 114093 3846 122439 3848
rect 114093 3843 114159 3846
rect 122373 3843 122439 3846
rect 80605 3770 80671 3773
rect 160185 3770 160251 3773
rect 80605 3768 160251 3770
rect 80605 3712 80610 3768
rect 80666 3712 160190 3768
rect 160246 3712 160251 3768
rect 80605 3710 160251 3712
rect 80605 3707 80671 3710
rect 160185 3707 160251 3710
rect 106181 3634 106247 3637
rect 426157 3634 426223 3637
rect 106181 3632 426223 3634
rect 106181 3576 106186 3632
rect 106242 3576 426162 3632
rect 426218 3576 426223 3632
rect 106181 3574 426223 3576
rect 106181 3571 106247 3574
rect 426157 3571 426223 3574
rect 110689 3498 110755 3501
rect 454493 3498 454559 3501
rect 110689 3496 454559 3498
rect 110689 3440 110694 3496
rect 110750 3440 454498 3496
rect 454554 3440 454559 3496
rect 110689 3438 454559 3440
rect 110689 3435 110755 3438
rect 454493 3435 454559 3438
rect 99557 3362 99623 3365
rect 109033 3362 109099 3365
rect 99557 3360 109099 3362
rect 99557 3304 99562 3360
rect 99618 3304 109038 3360
rect 109094 3304 109099 3360
rect 99557 3302 109099 3304
rect 99557 3299 99623 3302
rect 109033 3299 109099 3302
rect 111701 3362 111767 3365
rect 461577 3362 461643 3365
rect 111701 3360 461643 3362
rect 111701 3304 111706 3360
rect 111762 3304 461582 3360
rect 461638 3304 461643 3360
rect 111701 3302 461643 3304
rect 111701 3299 111767 3302
rect 461577 3299 461643 3302
rect 104433 3226 104499 3229
rect 111793 3226 111859 3229
rect 104433 3224 111859 3226
rect 104433 3168 104438 3224
rect 104494 3168 111798 3224
rect 111854 3168 111859 3224
rect 104433 3166 111859 3168
rect 104433 3163 104499 3166
rect 111793 3163 111859 3166
rect 95233 2818 95299 2821
rect 112621 2818 112687 2821
rect 95233 2816 100770 2818
rect 95233 2760 95238 2816
rect 95294 2760 100770 2816
rect 95233 2758 100770 2760
rect 95233 2755 95299 2758
rect 100710 2682 100770 2758
rect 108024 2816 112687 2818
rect 108024 2760 112626 2816
rect 112682 2760 112687 2816
rect 108024 2758 112687 2760
rect 108024 2682 108084 2758
rect 112621 2755 112687 2758
rect 100710 2622 108084 2682
rect 109033 2682 109099 2685
rect 115841 2682 115907 2685
rect 109033 2680 115907 2682
rect 109033 2624 109038 2680
rect 109094 2624 115846 2680
rect 115902 2624 115907 2680
rect 109033 2622 115907 2624
rect 109033 2619 109099 2622
rect 115841 2619 115907 2622
rect 127065 2682 127131 2685
rect 552565 2682 552631 2685
rect 127065 2680 552631 2682
rect 127065 2624 127070 2680
rect 127126 2624 552570 2680
rect 552626 2624 552631 2680
rect 127065 2622 552631 2624
rect 127065 2619 127131 2622
rect 552565 2619 552631 2622
rect 86677 2546 86743 2549
rect 104249 2546 104315 2549
rect 86677 2544 104315 2546
rect 86677 2488 86682 2544
rect 86738 2488 104254 2544
rect 104310 2488 104315 2544
rect 86677 2486 104315 2488
rect 86677 2483 86743 2486
rect 104249 2483 104315 2486
rect 107653 2546 107719 2549
rect 117957 2546 118023 2549
rect 107653 2544 118023 2546
rect 107653 2488 107658 2544
rect 107714 2488 117962 2544
rect 118018 2488 118023 2544
rect 107653 2486 118023 2488
rect 107653 2483 107719 2486
rect 117957 2483 118023 2486
rect 118141 2546 118207 2549
rect 146569 2546 146635 2549
rect 118141 2544 146635 2546
rect 118141 2488 118146 2544
rect 118202 2488 146574 2544
rect 146630 2488 146635 2544
rect 118141 2486 146635 2488
rect 118141 2483 118207 2486
rect 146569 2483 146635 2486
rect 56501 2410 56567 2413
rect 122097 2410 122163 2413
rect 56501 2408 122163 2410
rect 56501 2352 56506 2408
rect 56562 2352 122102 2408
rect 122158 2352 122163 2408
rect 56501 2350 122163 2352
rect 56501 2347 56567 2350
rect 122097 2347 122163 2350
rect 123569 2410 123635 2413
rect 145005 2410 145071 2413
rect 123569 2408 145071 2410
rect 123569 2352 123574 2408
rect 123630 2352 145010 2408
rect 145066 2352 145071 2408
rect 123569 2350 145071 2352
rect 123569 2347 123635 2350
rect 145005 2347 145071 2350
rect 110413 2274 110479 2277
rect 113357 2274 113423 2277
rect 110413 2272 113423 2274
rect 110413 2216 110418 2272
rect 110474 2216 113362 2272
rect 113418 2216 113423 2272
rect 110413 2214 113423 2216
rect 110413 2211 110479 2214
rect 113357 2211 113423 2214
rect 93117 2138 93183 2141
rect 299657 2138 299723 2141
rect 93117 2136 299723 2138
rect 93117 2080 93122 2136
rect 93178 2080 299662 2136
rect 299718 2080 299723 2136
rect 93117 2078 299723 2080
rect 93117 2075 93183 2078
rect 299657 2075 299723 2078
rect 100385 2002 100451 2005
rect 335077 2002 335143 2005
rect 100385 2000 335143 2002
rect 100385 1944 100390 2000
rect 100446 1944 335082 2000
rect 335138 1944 335143 2000
rect 100385 1942 335143 1944
rect 100385 1939 100451 1942
rect 335077 1939 335143 1942
rect 124121 1594 124187 1597
rect 126973 1594 127039 1597
rect 124121 1592 127039 1594
rect 124121 1536 124126 1592
rect 124182 1536 126978 1592
rect 127034 1536 127039 1592
rect 124121 1534 127039 1536
rect 124121 1531 124187 1534
rect 126973 1531 127039 1534
rect 111793 1322 111859 1325
rect 122833 1322 122899 1325
rect 111793 1320 122899 1322
rect 111793 1264 111798 1320
rect 111854 1264 122838 1320
rect 122894 1264 122899 1320
rect 111793 1262 122899 1264
rect 111793 1259 111859 1262
rect 122833 1259 122899 1262
rect 129641 1322 129707 1325
rect 136541 1322 136607 1325
rect 129641 1320 136607 1322
rect 129641 1264 129646 1320
rect 129702 1264 136546 1320
rect 136602 1264 136607 1320
rect 129641 1262 136607 1264
rect 129641 1259 129707 1262
rect 136541 1259 136607 1262
rect 89805 1186 89871 1189
rect 313273 1186 313339 1189
rect 89805 1184 313339 1186
rect 89805 1128 89810 1184
rect 89866 1128 313278 1184
rect 313334 1128 313339 1184
rect 89805 1126 313339 1128
rect 89805 1123 89871 1126
rect 313273 1123 313339 1126
rect 105261 1050 105327 1053
rect 135069 1050 135135 1053
rect 105261 1048 135135 1050
rect 105261 992 105266 1048
rect 105322 992 135074 1048
rect 135130 992 135135 1048
rect 105261 990 135135 992
rect 105261 987 105327 990
rect 135069 987 135135 990
rect 99741 914 99807 917
rect 384389 914 384455 917
rect 99741 912 384455 914
rect 99741 856 99746 912
rect 99802 856 384394 912
rect 384450 856 384455 912
rect 99741 854 384455 856
rect 99741 851 99807 854
rect 384389 851 384455 854
rect 93669 234 93735 237
rect 345381 234 345447 237
rect 93669 232 345447 234
rect 93669 176 93674 232
rect 93730 176 345386 232
rect 345442 176 345447 232
rect 93669 174 345447 176
rect 93669 171 93735 174
rect 345381 171 345447 174
rect 126421 98 126487 101
rect 556337 98 556403 101
rect 126421 96 556403 98
rect 126421 40 126426 96
rect 126482 40 556342 96
rect 556398 40 556403 96
rect 126421 38 556403 40
rect 126421 35 126487 38
rect 556337 35 556403 38
<< via3 >>
rect 31892 154396 31956 154460
rect 25820 153580 25884 153644
rect 143580 153172 143644 153236
rect 139348 152900 139412 152964
rect 37596 152356 37660 152420
rect 137876 152492 137940 152556
rect 19932 152084 19996 152148
rect 37596 151948 37660 152012
rect 35756 151812 35820 151876
rect 136588 151812 136652 151876
rect 25820 151676 25884 151740
rect 143580 151676 143644 151740
rect 31892 151540 31956 151604
rect 136588 151540 136652 151604
rect 35756 151404 35820 151468
rect 139348 151404 139412 151468
rect 137876 151268 137940 151332
rect 151124 24924 151188 24988
rect 151124 17716 151188 17780
rect 19932 14588 19996 14652
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 154746 20414 164898
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 154746 24914 169398
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 154746 29414 173898
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 154746 33914 178398
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 154746 38414 182898
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 154746 42914 187398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 154746 47414 155898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 154746 51914 160398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 154746 56414 164898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 154746 60914 169398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 154746 65414 173898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 154746 69914 178398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 154746 74414 182898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 154746 78914 187398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 154746 83414 155898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 154746 87914 160398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 154746 92414 164898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 154746 96914 169398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 154746 101414 173898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 154746 105914 178398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 154746 110414 182898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 154746 114914 187398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 154746 119414 155898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 154746 123914 160398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 154746 128414 164898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 154746 132914 169398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 154746 137414 173898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 154746 141914 178398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 154746 146414 182898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 154746 150914 187398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 31891 154460 31957 154461
rect 31891 154396 31892 154460
rect 31956 154396 31957 154460
rect 31891 154395 31957 154396
rect 25819 153644 25885 153645
rect 25819 153580 25820 153644
rect 25884 153580 25885 153644
rect 25819 153579 25885 153580
rect 19931 152148 19997 152149
rect 19931 152084 19932 152148
rect 19996 152084 19997 152148
rect 19931 152083 19997 152084
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 19934 14653 19994 152083
rect 25822 151741 25882 153579
rect 25819 151740 25885 151741
rect 25819 151676 25820 151740
rect 25884 151676 25885 151740
rect 25819 151675 25885 151676
rect 31894 151605 31954 154395
rect 143579 153236 143645 153237
rect 143579 153172 143580 153236
rect 143644 153172 143645 153236
rect 143579 153171 143645 153172
rect 139347 152964 139413 152965
rect 139347 152900 139348 152964
rect 139412 152900 139413 152964
rect 139347 152899 139413 152900
rect 137875 152556 137941 152557
rect 137875 152492 137876 152556
rect 137940 152492 137941 152556
rect 137875 152491 137941 152492
rect 37595 152420 37661 152421
rect 37595 152356 37596 152420
rect 37660 152356 37661 152420
rect 37595 152355 37661 152356
rect 37598 152013 37658 152355
rect 37595 152012 37661 152013
rect 37595 151948 37596 152012
rect 37660 151948 37661 152012
rect 37595 151947 37661 151948
rect 35755 151876 35821 151877
rect 35755 151812 35756 151876
rect 35820 151812 35821 151876
rect 35755 151811 35821 151812
rect 136587 151876 136653 151877
rect 136587 151812 136588 151876
rect 136652 151812 136653 151876
rect 136587 151811 136653 151812
rect 31891 151604 31957 151605
rect 31891 151540 31892 151604
rect 31956 151540 31957 151604
rect 31891 151539 31957 151540
rect 35758 151469 35818 151811
rect 136590 151605 136650 151811
rect 136587 151604 136653 151605
rect 136587 151540 136588 151604
rect 136652 151540 136653 151604
rect 136587 151539 136653 151540
rect 35755 151468 35821 151469
rect 35755 151404 35756 151468
rect 35820 151404 35821 151468
rect 35755 151403 35821 151404
rect 137878 151333 137938 152491
rect 139350 151469 139410 152899
rect 143582 151741 143642 153171
rect 143579 151740 143645 151741
rect 143579 151676 143580 151740
rect 143644 151676 143645 151740
rect 143579 151675 143645 151676
rect 139347 151468 139413 151469
rect 139347 151404 139348 151468
rect 139412 151404 139413 151468
rect 139347 151403 139413 151404
rect 137875 151332 137941 151333
rect 137875 151268 137876 151332
rect 137940 151268 137941 151332
rect 137875 151267 137941 151268
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 39568 115954 39888 115986
rect 39568 115718 39610 115954
rect 39846 115718 39888 115954
rect 39568 115634 39888 115718
rect 39568 115398 39610 115634
rect 39846 115398 39888 115634
rect 39568 115366 39888 115398
rect 70288 115954 70608 115986
rect 70288 115718 70330 115954
rect 70566 115718 70608 115954
rect 70288 115634 70608 115718
rect 70288 115398 70330 115634
rect 70566 115398 70608 115634
rect 70288 115366 70608 115398
rect 101008 115954 101328 115986
rect 101008 115718 101050 115954
rect 101286 115718 101328 115954
rect 101008 115634 101328 115718
rect 101008 115398 101050 115634
rect 101286 115398 101328 115634
rect 101008 115366 101328 115398
rect 131728 115954 132048 115986
rect 131728 115718 131770 115954
rect 132006 115718 132048 115954
rect 131728 115634 132048 115718
rect 131728 115398 131770 115634
rect 132006 115398 132048 115634
rect 131728 115366 132048 115398
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 39568 79954 39888 79986
rect 39568 79718 39610 79954
rect 39846 79718 39888 79954
rect 39568 79634 39888 79718
rect 39568 79398 39610 79634
rect 39846 79398 39888 79634
rect 39568 79366 39888 79398
rect 70288 79954 70608 79986
rect 70288 79718 70330 79954
rect 70566 79718 70608 79954
rect 70288 79634 70608 79718
rect 70288 79398 70330 79634
rect 70566 79398 70608 79634
rect 70288 79366 70608 79398
rect 101008 79954 101328 79986
rect 101008 79718 101050 79954
rect 101286 79718 101328 79954
rect 101008 79634 101328 79718
rect 101008 79398 101050 79634
rect 101286 79398 101328 79634
rect 101008 79366 101328 79398
rect 131728 79954 132048 79986
rect 131728 79718 131770 79954
rect 132006 79718 132048 79954
rect 131728 79634 132048 79718
rect 131728 79398 131770 79634
rect 132006 79398 132048 79634
rect 131728 79366 132048 79398
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 39568 43954 39888 43986
rect 39568 43718 39610 43954
rect 39846 43718 39888 43954
rect 39568 43634 39888 43718
rect 39568 43398 39610 43634
rect 39846 43398 39888 43634
rect 39568 43366 39888 43398
rect 70288 43954 70608 43986
rect 70288 43718 70330 43954
rect 70566 43718 70608 43954
rect 70288 43634 70608 43718
rect 70288 43398 70330 43634
rect 70566 43398 70608 43634
rect 70288 43366 70608 43398
rect 101008 43954 101328 43986
rect 101008 43718 101050 43954
rect 101286 43718 101328 43954
rect 101008 43634 101328 43718
rect 101008 43398 101050 43634
rect 101286 43398 101328 43634
rect 101008 43366 101328 43398
rect 131728 43954 132048 43986
rect 131728 43718 131770 43954
rect 132006 43718 132048 43954
rect 131728 43634 132048 43718
rect 131728 43398 131770 43634
rect 132006 43398 132048 43634
rect 131728 43366 132048 43398
rect 24208 39454 24528 39486
rect 24208 39218 24250 39454
rect 24486 39218 24528 39454
rect 24208 39134 24528 39218
rect 24208 38898 24250 39134
rect 24486 38898 24528 39134
rect 24208 38866 24528 38898
rect 54928 39454 55248 39486
rect 54928 39218 54970 39454
rect 55206 39218 55248 39454
rect 54928 39134 55248 39218
rect 54928 38898 54970 39134
rect 55206 38898 55248 39134
rect 54928 38866 55248 38898
rect 85648 39454 85968 39486
rect 85648 39218 85690 39454
rect 85926 39218 85968 39454
rect 85648 39134 85968 39218
rect 85648 38898 85690 39134
rect 85926 38898 85968 39134
rect 85648 38866 85968 38898
rect 116368 39454 116688 39486
rect 116368 39218 116410 39454
rect 116646 39218 116688 39454
rect 116368 39134 116688 39218
rect 116368 38898 116410 39134
rect 116646 38898 116688 39134
rect 116368 38866 116688 38898
rect 147088 39454 147408 39486
rect 147088 39218 147130 39454
rect 147366 39218 147408 39454
rect 147088 39134 147408 39218
rect 147088 38898 147130 39134
rect 147366 38898 147408 39134
rect 147088 38866 147408 38898
rect 151123 24988 151189 24989
rect 151123 24924 151124 24988
rect 151188 24924 151189 24988
rect 151123 24923 151189 24924
rect 19931 14652 19997 14653
rect 19931 14588 19932 14652
rect 19996 14588 19997 14652
rect 19931 14587 19997 14588
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 37794 3454 38414 18000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 7954 42914 18000
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 12454 47414 18000
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 16954 51914 18000
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 73794 3454 74414 18000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 7954 78914 18000
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 12454 83414 18000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 16954 87914 18000
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 109794 3454 110414 18000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 7954 114914 18000
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 18000
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 16954 123914 18000
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 145794 3454 146414 18000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 18000
rect 151126 17781 151186 24923
rect 151123 17780 151189 17781
rect 151123 17716 151124 17780
rect 151188 17716 151189 17780
rect 151123 17715 151189 17716
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 39610 115718 39846 115954
rect 39610 115398 39846 115634
rect 70330 115718 70566 115954
rect 70330 115398 70566 115634
rect 101050 115718 101286 115954
rect 101050 115398 101286 115634
rect 131770 115718 132006 115954
rect 131770 115398 132006 115634
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 39610 79718 39846 79954
rect 39610 79398 39846 79634
rect 70330 79718 70566 79954
rect 70330 79398 70566 79634
rect 101050 79718 101286 79954
rect 101050 79398 101286 79634
rect 131770 79718 132006 79954
rect 131770 79398 132006 79634
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 39610 43718 39846 43954
rect 39610 43398 39846 43634
rect 70330 43718 70566 43954
rect 70330 43398 70566 43634
rect 101050 43718 101286 43954
rect 101050 43398 101286 43634
rect 131770 43718 132006 43954
rect 131770 43398 132006 43634
rect 24250 39218 24486 39454
rect 24250 38898 24486 39134
rect 54970 39218 55206 39454
rect 54970 38898 55206 39134
rect 85690 39218 85926 39454
rect 85690 38898 85926 39134
rect 116410 39218 116646 39454
rect 116410 38898 116646 39134
rect 147130 39218 147366 39454
rect 147130 38898 147366 39134
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 39610 115954
rect 39846 115718 70330 115954
rect 70566 115718 101050 115954
rect 101286 115718 131770 115954
rect 132006 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 39610 115634
rect 39846 115398 70330 115634
rect 70566 115398 101050 115634
rect 101286 115398 131770 115634
rect 132006 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 39610 79954
rect 39846 79718 70330 79954
rect 70566 79718 101050 79954
rect 101286 79718 131770 79954
rect 132006 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 39610 79634
rect 39846 79398 70330 79634
rect 70566 79398 101050 79634
rect 101286 79398 131770 79634
rect 132006 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 39610 43954
rect 39846 43718 70330 43954
rect 70566 43718 101050 43954
rect 101286 43718 131770 43954
rect 132006 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 39610 43634
rect 39846 43398 70330 43634
rect 70566 43398 101050 43634
rect 101286 43398 131770 43634
rect 132006 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 24250 39454
rect 24486 39218 54970 39454
rect 55206 39218 85690 39454
rect 85926 39218 116410 39454
rect 116646 39218 147130 39454
rect 147366 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 24250 39134
rect 24486 38898 54970 39134
rect 55206 38898 85690 39134
rect 85926 38898 116410 39134
rect 116646 38898 147130 39134
rect 147366 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sha1_top  sha1_top_inst
timestamp 0
transform 1 0 20000 0 1 20000
box 238 0 130608 132746
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 18000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 154746 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 18000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 154746 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 18000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 154746 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 18000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 154746 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 18000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 154746 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 18000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 154746 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 18000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 154746 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 154746 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 154746 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 154746 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 154746 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 154746 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 154746 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 154746 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 154746 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 154746 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 154746 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 154746 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 154746 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 154746 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 154746 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 154746 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 154746 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 18000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 154746 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 18000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 154746 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 18000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 154746 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 18000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 154746 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 18000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 154746 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 18000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 154746 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 18000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 154746 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
