magic
tech sky130A
magscale 1 2
timestamp 1652849600
<< obsli1 >>
rect 1104 2159 91540 92497
<< obsm1 >>
rect 106 8 92538 92528
<< metal2 >>
rect 386 94000 442 94800
rect 1122 94000 1178 94800
rect 1950 94000 2006 94800
rect 2778 94000 2834 94800
rect 3606 94000 3662 94800
rect 4434 94000 4490 94800
rect 5262 94000 5318 94800
rect 5998 94000 6054 94800
rect 6826 94000 6882 94800
rect 7654 94000 7710 94800
rect 8482 94000 8538 94800
rect 9310 94000 9366 94800
rect 10138 94000 10194 94800
rect 10874 94000 10930 94800
rect 11702 94000 11758 94800
rect 12530 94000 12586 94800
rect 13358 94000 13414 94800
rect 14186 94000 14242 94800
rect 15014 94000 15070 94800
rect 15750 94000 15806 94800
rect 16578 94000 16634 94800
rect 17406 94000 17462 94800
rect 18234 94000 18290 94800
rect 19062 94000 19118 94800
rect 19890 94000 19946 94800
rect 20626 94000 20682 94800
rect 21454 94000 21510 94800
rect 22282 94000 22338 94800
rect 23110 94000 23166 94800
rect 23938 94000 23994 94800
rect 24766 94000 24822 94800
rect 25502 94000 25558 94800
rect 26330 94000 26386 94800
rect 27158 94000 27214 94800
rect 27986 94000 28042 94800
rect 28814 94000 28870 94800
rect 29642 94000 29698 94800
rect 30378 94000 30434 94800
rect 31206 94000 31262 94800
rect 32034 94000 32090 94800
rect 32862 94000 32918 94800
rect 33690 94000 33746 94800
rect 34518 94000 34574 94800
rect 35254 94000 35310 94800
rect 36082 94000 36138 94800
rect 36910 94000 36966 94800
rect 37738 94000 37794 94800
rect 38566 94000 38622 94800
rect 39394 94000 39450 94800
rect 40130 94000 40186 94800
rect 40958 94000 41014 94800
rect 41786 94000 41842 94800
rect 42614 94000 42670 94800
rect 43442 94000 43498 94800
rect 44270 94000 44326 94800
rect 45006 94000 45062 94800
rect 45834 94000 45890 94800
rect 46662 94000 46718 94800
rect 47490 94000 47546 94800
rect 48318 94000 48374 94800
rect 49146 94000 49202 94800
rect 49882 94000 49938 94800
rect 50710 94000 50766 94800
rect 51538 94000 51594 94800
rect 52366 94000 52422 94800
rect 53194 94000 53250 94800
rect 54022 94000 54078 94800
rect 54758 94000 54814 94800
rect 55586 94000 55642 94800
rect 56414 94000 56470 94800
rect 57242 94000 57298 94800
rect 58070 94000 58126 94800
rect 58898 94000 58954 94800
rect 59634 94000 59690 94800
rect 60462 94000 60518 94800
rect 61290 94000 61346 94800
rect 62118 94000 62174 94800
rect 62946 94000 63002 94800
rect 63774 94000 63830 94800
rect 64510 94000 64566 94800
rect 65338 94000 65394 94800
rect 66166 94000 66222 94800
rect 66994 94000 67050 94800
rect 67822 94000 67878 94800
rect 68650 94000 68706 94800
rect 69386 94000 69442 94800
rect 70214 94000 70270 94800
rect 71042 94000 71098 94800
rect 71870 94000 71926 94800
rect 72698 94000 72754 94800
rect 73526 94000 73582 94800
rect 74262 94000 74318 94800
rect 75090 94000 75146 94800
rect 75918 94000 75974 94800
rect 76746 94000 76802 94800
rect 77574 94000 77630 94800
rect 78402 94000 78458 94800
rect 79138 94000 79194 94800
rect 79966 94000 80022 94800
rect 80794 94000 80850 94800
rect 81622 94000 81678 94800
rect 82450 94000 82506 94800
rect 83278 94000 83334 94800
rect 84014 94000 84070 94800
rect 84842 94000 84898 94800
rect 85670 94000 85726 94800
rect 86498 94000 86554 94800
rect 87326 94000 87382 94800
rect 88154 94000 88210 94800
rect 88890 94000 88946 94800
rect 89718 94000 89774 94800
rect 90546 94000 90602 94800
rect 91374 94000 91430 94800
rect 92202 94000 92258 94800
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68282 0 68338 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77850 0 77906 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78402 0 78458 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87418 0 87474 800
rect 87602 0 87658 800
rect 87786 0 87842 800
rect 87970 0 88026 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90638 0 90694 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92478 0 92534 800
<< obsm2 >>
rect 112 93944 330 94058
rect 498 93944 1066 94058
rect 1234 93944 1894 94058
rect 2062 93944 2722 94058
rect 2890 93944 3550 94058
rect 3718 93944 4378 94058
rect 4546 93944 5206 94058
rect 5374 93944 5942 94058
rect 6110 93944 6770 94058
rect 6938 93944 7598 94058
rect 7766 93944 8426 94058
rect 8594 93944 9254 94058
rect 9422 93944 10082 94058
rect 10250 93944 10818 94058
rect 10986 93944 11646 94058
rect 11814 93944 12474 94058
rect 12642 93944 13302 94058
rect 13470 93944 14130 94058
rect 14298 93944 14958 94058
rect 15126 93944 15694 94058
rect 15862 93944 16522 94058
rect 16690 93944 17350 94058
rect 17518 93944 18178 94058
rect 18346 93944 19006 94058
rect 19174 93944 19834 94058
rect 20002 93944 20570 94058
rect 20738 93944 21398 94058
rect 21566 93944 22226 94058
rect 22394 93944 23054 94058
rect 23222 93944 23882 94058
rect 24050 93944 24710 94058
rect 24878 93944 25446 94058
rect 25614 93944 26274 94058
rect 26442 93944 27102 94058
rect 27270 93944 27930 94058
rect 28098 93944 28758 94058
rect 28926 93944 29586 94058
rect 29754 93944 30322 94058
rect 30490 93944 31150 94058
rect 31318 93944 31978 94058
rect 32146 93944 32806 94058
rect 32974 93944 33634 94058
rect 33802 93944 34462 94058
rect 34630 93944 35198 94058
rect 35366 93944 36026 94058
rect 36194 93944 36854 94058
rect 37022 93944 37682 94058
rect 37850 93944 38510 94058
rect 38678 93944 39338 94058
rect 39506 93944 40074 94058
rect 40242 93944 40902 94058
rect 41070 93944 41730 94058
rect 41898 93944 42558 94058
rect 42726 93944 43386 94058
rect 43554 93944 44214 94058
rect 44382 93944 44950 94058
rect 45118 93944 45778 94058
rect 45946 93944 46606 94058
rect 46774 93944 47434 94058
rect 47602 93944 48262 94058
rect 48430 93944 49090 94058
rect 49258 93944 49826 94058
rect 49994 93944 50654 94058
rect 50822 93944 51482 94058
rect 51650 93944 52310 94058
rect 52478 93944 53138 94058
rect 53306 93944 53966 94058
rect 54134 93944 54702 94058
rect 54870 93944 55530 94058
rect 55698 93944 56358 94058
rect 56526 93944 57186 94058
rect 57354 93944 58014 94058
rect 58182 93944 58842 94058
rect 59010 93944 59578 94058
rect 59746 93944 60406 94058
rect 60574 93944 61234 94058
rect 61402 93944 62062 94058
rect 62230 93944 62890 94058
rect 63058 93944 63718 94058
rect 63886 93944 64454 94058
rect 64622 93944 65282 94058
rect 65450 93944 66110 94058
rect 66278 93944 66938 94058
rect 67106 93944 67766 94058
rect 67934 93944 68594 94058
rect 68762 93944 69330 94058
rect 69498 93944 70158 94058
rect 70326 93944 70986 94058
rect 71154 93944 71814 94058
rect 71982 93944 72642 94058
rect 72810 93944 73470 94058
rect 73638 93944 74206 94058
rect 74374 93944 75034 94058
rect 75202 93944 75862 94058
rect 76030 93944 76690 94058
rect 76858 93944 77518 94058
rect 77686 93944 78346 94058
rect 78514 93944 79082 94058
rect 79250 93944 79910 94058
rect 80078 93944 80738 94058
rect 80906 93944 81566 94058
rect 81734 93944 82394 94058
rect 82562 93944 83222 94058
rect 83390 93944 83958 94058
rect 84126 93944 84786 94058
rect 84954 93944 85614 94058
rect 85782 93944 86442 94058
rect 86610 93944 87270 94058
rect 87438 93944 88098 94058
rect 88266 93944 88834 94058
rect 89002 93944 89662 94058
rect 89830 93944 90490 94058
rect 90658 93944 91318 94058
rect 91486 93944 92146 94058
rect 92314 93944 92532 94058
rect 112 856 92532 93944
rect 222 2 238 856
rect 406 2 422 856
rect 590 2 606 856
rect 774 2 790 856
rect 958 2 974 856
rect 1142 2 1158 856
rect 1326 2 1342 856
rect 1510 2 1526 856
rect 1694 2 1710 856
rect 1878 2 1894 856
rect 2062 2 2078 856
rect 2246 2 2262 856
rect 2430 2 2446 856
rect 2614 2 2630 856
rect 2798 2 2814 856
rect 2982 2 2998 856
rect 3166 2 3182 856
rect 3350 2 3366 856
rect 3534 2 3550 856
rect 3718 2 3734 856
rect 3902 2 3918 856
rect 4086 2 4102 856
rect 4270 2 4286 856
rect 4454 2 4562 856
rect 4730 2 4746 856
rect 4914 2 4930 856
rect 5098 2 5114 856
rect 5282 2 5298 856
rect 5466 2 5482 856
rect 5650 2 5666 856
rect 5834 2 5850 856
rect 6018 2 6034 856
rect 6202 2 6218 856
rect 6386 2 6402 856
rect 6570 2 6586 856
rect 6754 2 6770 856
rect 6938 2 6954 856
rect 7122 2 7138 856
rect 7306 2 7322 856
rect 7490 2 7506 856
rect 7674 2 7690 856
rect 7858 2 7874 856
rect 8042 2 8058 856
rect 8226 2 8242 856
rect 8410 2 8426 856
rect 8594 2 8610 856
rect 8778 2 8886 856
rect 9054 2 9070 856
rect 9238 2 9254 856
rect 9422 2 9438 856
rect 9606 2 9622 856
rect 9790 2 9806 856
rect 9974 2 9990 856
rect 10158 2 10174 856
rect 10342 2 10358 856
rect 10526 2 10542 856
rect 10710 2 10726 856
rect 10894 2 10910 856
rect 11078 2 11094 856
rect 11262 2 11278 856
rect 11446 2 11462 856
rect 11630 2 11646 856
rect 11814 2 11830 856
rect 11998 2 12014 856
rect 12182 2 12198 856
rect 12366 2 12382 856
rect 12550 2 12566 856
rect 12734 2 12750 856
rect 12918 2 12934 856
rect 13102 2 13118 856
rect 13286 2 13394 856
rect 13562 2 13578 856
rect 13746 2 13762 856
rect 13930 2 13946 856
rect 14114 2 14130 856
rect 14298 2 14314 856
rect 14482 2 14498 856
rect 14666 2 14682 856
rect 14850 2 14866 856
rect 15034 2 15050 856
rect 15218 2 15234 856
rect 15402 2 15418 856
rect 15586 2 15602 856
rect 15770 2 15786 856
rect 15954 2 15970 856
rect 16138 2 16154 856
rect 16322 2 16338 856
rect 16506 2 16522 856
rect 16690 2 16706 856
rect 16874 2 16890 856
rect 17058 2 17074 856
rect 17242 2 17258 856
rect 17426 2 17442 856
rect 17610 2 17718 856
rect 17886 2 17902 856
rect 18070 2 18086 856
rect 18254 2 18270 856
rect 18438 2 18454 856
rect 18622 2 18638 856
rect 18806 2 18822 856
rect 18990 2 19006 856
rect 19174 2 19190 856
rect 19358 2 19374 856
rect 19542 2 19558 856
rect 19726 2 19742 856
rect 19910 2 19926 856
rect 20094 2 20110 856
rect 20278 2 20294 856
rect 20462 2 20478 856
rect 20646 2 20662 856
rect 20830 2 20846 856
rect 21014 2 21030 856
rect 21198 2 21214 856
rect 21382 2 21398 856
rect 21566 2 21582 856
rect 21750 2 21766 856
rect 21934 2 21950 856
rect 22118 2 22226 856
rect 22394 2 22410 856
rect 22578 2 22594 856
rect 22762 2 22778 856
rect 22946 2 22962 856
rect 23130 2 23146 856
rect 23314 2 23330 856
rect 23498 2 23514 856
rect 23682 2 23698 856
rect 23866 2 23882 856
rect 24050 2 24066 856
rect 24234 2 24250 856
rect 24418 2 24434 856
rect 24602 2 24618 856
rect 24786 2 24802 856
rect 24970 2 24986 856
rect 25154 2 25170 856
rect 25338 2 25354 856
rect 25522 2 25538 856
rect 25706 2 25722 856
rect 25890 2 25906 856
rect 26074 2 26090 856
rect 26258 2 26274 856
rect 26442 2 26550 856
rect 26718 2 26734 856
rect 26902 2 26918 856
rect 27086 2 27102 856
rect 27270 2 27286 856
rect 27454 2 27470 856
rect 27638 2 27654 856
rect 27822 2 27838 856
rect 28006 2 28022 856
rect 28190 2 28206 856
rect 28374 2 28390 856
rect 28558 2 28574 856
rect 28742 2 28758 856
rect 28926 2 28942 856
rect 29110 2 29126 856
rect 29294 2 29310 856
rect 29478 2 29494 856
rect 29662 2 29678 856
rect 29846 2 29862 856
rect 30030 2 30046 856
rect 30214 2 30230 856
rect 30398 2 30414 856
rect 30582 2 30598 856
rect 30766 2 30782 856
rect 30950 2 31058 856
rect 31226 2 31242 856
rect 31410 2 31426 856
rect 31594 2 31610 856
rect 31778 2 31794 856
rect 31962 2 31978 856
rect 32146 2 32162 856
rect 32330 2 32346 856
rect 32514 2 32530 856
rect 32698 2 32714 856
rect 32882 2 32898 856
rect 33066 2 33082 856
rect 33250 2 33266 856
rect 33434 2 33450 856
rect 33618 2 33634 856
rect 33802 2 33818 856
rect 33986 2 34002 856
rect 34170 2 34186 856
rect 34354 2 34370 856
rect 34538 2 34554 856
rect 34722 2 34738 856
rect 34906 2 34922 856
rect 35090 2 35106 856
rect 35274 2 35382 856
rect 35550 2 35566 856
rect 35734 2 35750 856
rect 35918 2 35934 856
rect 36102 2 36118 856
rect 36286 2 36302 856
rect 36470 2 36486 856
rect 36654 2 36670 856
rect 36838 2 36854 856
rect 37022 2 37038 856
rect 37206 2 37222 856
rect 37390 2 37406 856
rect 37574 2 37590 856
rect 37758 2 37774 856
rect 37942 2 37958 856
rect 38126 2 38142 856
rect 38310 2 38326 856
rect 38494 2 38510 856
rect 38678 2 38694 856
rect 38862 2 38878 856
rect 39046 2 39062 856
rect 39230 2 39246 856
rect 39414 2 39430 856
rect 39598 2 39614 856
rect 39782 2 39890 856
rect 40058 2 40074 856
rect 40242 2 40258 856
rect 40426 2 40442 856
rect 40610 2 40626 856
rect 40794 2 40810 856
rect 40978 2 40994 856
rect 41162 2 41178 856
rect 41346 2 41362 856
rect 41530 2 41546 856
rect 41714 2 41730 856
rect 41898 2 41914 856
rect 42082 2 42098 856
rect 42266 2 42282 856
rect 42450 2 42466 856
rect 42634 2 42650 856
rect 42818 2 42834 856
rect 43002 2 43018 856
rect 43186 2 43202 856
rect 43370 2 43386 856
rect 43554 2 43570 856
rect 43738 2 43754 856
rect 43922 2 43938 856
rect 44106 2 44214 856
rect 44382 2 44398 856
rect 44566 2 44582 856
rect 44750 2 44766 856
rect 44934 2 44950 856
rect 45118 2 45134 856
rect 45302 2 45318 856
rect 45486 2 45502 856
rect 45670 2 45686 856
rect 45854 2 45870 856
rect 46038 2 46054 856
rect 46222 2 46238 856
rect 46406 2 46422 856
rect 46590 2 46606 856
rect 46774 2 46790 856
rect 46958 2 46974 856
rect 47142 2 47158 856
rect 47326 2 47342 856
rect 47510 2 47526 856
rect 47694 2 47710 856
rect 47878 2 47894 856
rect 48062 2 48078 856
rect 48246 2 48262 856
rect 48430 2 48446 856
rect 48614 2 48722 856
rect 48890 2 48906 856
rect 49074 2 49090 856
rect 49258 2 49274 856
rect 49442 2 49458 856
rect 49626 2 49642 856
rect 49810 2 49826 856
rect 49994 2 50010 856
rect 50178 2 50194 856
rect 50362 2 50378 856
rect 50546 2 50562 856
rect 50730 2 50746 856
rect 50914 2 50930 856
rect 51098 2 51114 856
rect 51282 2 51298 856
rect 51466 2 51482 856
rect 51650 2 51666 856
rect 51834 2 51850 856
rect 52018 2 52034 856
rect 52202 2 52218 856
rect 52386 2 52402 856
rect 52570 2 52586 856
rect 52754 2 52770 856
rect 52938 2 53046 856
rect 53214 2 53230 856
rect 53398 2 53414 856
rect 53582 2 53598 856
rect 53766 2 53782 856
rect 53950 2 53966 856
rect 54134 2 54150 856
rect 54318 2 54334 856
rect 54502 2 54518 856
rect 54686 2 54702 856
rect 54870 2 54886 856
rect 55054 2 55070 856
rect 55238 2 55254 856
rect 55422 2 55438 856
rect 55606 2 55622 856
rect 55790 2 55806 856
rect 55974 2 55990 856
rect 56158 2 56174 856
rect 56342 2 56358 856
rect 56526 2 56542 856
rect 56710 2 56726 856
rect 56894 2 56910 856
rect 57078 2 57094 856
rect 57262 2 57278 856
rect 57446 2 57554 856
rect 57722 2 57738 856
rect 57906 2 57922 856
rect 58090 2 58106 856
rect 58274 2 58290 856
rect 58458 2 58474 856
rect 58642 2 58658 856
rect 58826 2 58842 856
rect 59010 2 59026 856
rect 59194 2 59210 856
rect 59378 2 59394 856
rect 59562 2 59578 856
rect 59746 2 59762 856
rect 59930 2 59946 856
rect 60114 2 60130 856
rect 60298 2 60314 856
rect 60482 2 60498 856
rect 60666 2 60682 856
rect 60850 2 60866 856
rect 61034 2 61050 856
rect 61218 2 61234 856
rect 61402 2 61418 856
rect 61586 2 61602 856
rect 61770 2 61878 856
rect 62046 2 62062 856
rect 62230 2 62246 856
rect 62414 2 62430 856
rect 62598 2 62614 856
rect 62782 2 62798 856
rect 62966 2 62982 856
rect 63150 2 63166 856
rect 63334 2 63350 856
rect 63518 2 63534 856
rect 63702 2 63718 856
rect 63886 2 63902 856
rect 64070 2 64086 856
rect 64254 2 64270 856
rect 64438 2 64454 856
rect 64622 2 64638 856
rect 64806 2 64822 856
rect 64990 2 65006 856
rect 65174 2 65190 856
rect 65358 2 65374 856
rect 65542 2 65558 856
rect 65726 2 65742 856
rect 65910 2 65926 856
rect 66094 2 66110 856
rect 66278 2 66386 856
rect 66554 2 66570 856
rect 66738 2 66754 856
rect 66922 2 66938 856
rect 67106 2 67122 856
rect 67290 2 67306 856
rect 67474 2 67490 856
rect 67658 2 67674 856
rect 67842 2 67858 856
rect 68026 2 68042 856
rect 68210 2 68226 856
rect 68394 2 68410 856
rect 68578 2 68594 856
rect 68762 2 68778 856
rect 68946 2 68962 856
rect 69130 2 69146 856
rect 69314 2 69330 856
rect 69498 2 69514 856
rect 69682 2 69698 856
rect 69866 2 69882 856
rect 70050 2 70066 856
rect 70234 2 70250 856
rect 70418 2 70434 856
rect 70602 2 70710 856
rect 70878 2 70894 856
rect 71062 2 71078 856
rect 71246 2 71262 856
rect 71430 2 71446 856
rect 71614 2 71630 856
rect 71798 2 71814 856
rect 71982 2 71998 856
rect 72166 2 72182 856
rect 72350 2 72366 856
rect 72534 2 72550 856
rect 72718 2 72734 856
rect 72902 2 72918 856
rect 73086 2 73102 856
rect 73270 2 73286 856
rect 73454 2 73470 856
rect 73638 2 73654 856
rect 73822 2 73838 856
rect 74006 2 74022 856
rect 74190 2 74206 856
rect 74374 2 74390 856
rect 74558 2 74574 856
rect 74742 2 74758 856
rect 74926 2 74942 856
rect 75110 2 75218 856
rect 75386 2 75402 856
rect 75570 2 75586 856
rect 75754 2 75770 856
rect 75938 2 75954 856
rect 76122 2 76138 856
rect 76306 2 76322 856
rect 76490 2 76506 856
rect 76674 2 76690 856
rect 76858 2 76874 856
rect 77042 2 77058 856
rect 77226 2 77242 856
rect 77410 2 77426 856
rect 77594 2 77610 856
rect 77778 2 77794 856
rect 77962 2 77978 856
rect 78146 2 78162 856
rect 78330 2 78346 856
rect 78514 2 78530 856
rect 78698 2 78714 856
rect 78882 2 78898 856
rect 79066 2 79082 856
rect 79250 2 79266 856
rect 79434 2 79542 856
rect 79710 2 79726 856
rect 79894 2 79910 856
rect 80078 2 80094 856
rect 80262 2 80278 856
rect 80446 2 80462 856
rect 80630 2 80646 856
rect 80814 2 80830 856
rect 80998 2 81014 856
rect 81182 2 81198 856
rect 81366 2 81382 856
rect 81550 2 81566 856
rect 81734 2 81750 856
rect 81918 2 81934 856
rect 82102 2 82118 856
rect 82286 2 82302 856
rect 82470 2 82486 856
rect 82654 2 82670 856
rect 82838 2 82854 856
rect 83022 2 83038 856
rect 83206 2 83222 856
rect 83390 2 83406 856
rect 83574 2 83590 856
rect 83758 2 83774 856
rect 83942 2 84050 856
rect 84218 2 84234 856
rect 84402 2 84418 856
rect 84586 2 84602 856
rect 84770 2 84786 856
rect 84954 2 84970 856
rect 85138 2 85154 856
rect 85322 2 85338 856
rect 85506 2 85522 856
rect 85690 2 85706 856
rect 85874 2 85890 856
rect 86058 2 86074 856
rect 86242 2 86258 856
rect 86426 2 86442 856
rect 86610 2 86626 856
rect 86794 2 86810 856
rect 86978 2 86994 856
rect 87162 2 87178 856
rect 87346 2 87362 856
rect 87530 2 87546 856
rect 87714 2 87730 856
rect 87898 2 87914 856
rect 88082 2 88098 856
rect 88266 2 88374 856
rect 88542 2 88558 856
rect 88726 2 88742 856
rect 88910 2 88926 856
rect 89094 2 89110 856
rect 89278 2 89294 856
rect 89462 2 89478 856
rect 89646 2 89662 856
rect 89830 2 89846 856
rect 90014 2 90030 856
rect 90198 2 90214 856
rect 90382 2 90398 856
rect 90566 2 90582 856
rect 90750 2 90766 856
rect 90934 2 90950 856
rect 91118 2 91134 856
rect 91302 2 91318 856
rect 91486 2 91502 856
rect 91670 2 91686 856
rect 91854 2 91870 856
rect 92038 2 92054 856
rect 92222 2 92238 856
rect 92406 2 92422 856
<< obsm3 >>
rect 565 35 81328 92513
<< metal4 >>
rect 4208 2128 4528 92528
rect 19568 2128 19888 92528
rect 34928 2128 35248 92528
rect 50288 2128 50608 92528
rect 65648 2128 65968 92528
rect 81008 2128 81328 92528
<< obsm4 >>
rect 611 2048 4128 92173
rect 4608 2048 19488 92173
rect 19968 2048 34848 92173
rect 35328 2048 50208 92173
rect 50688 2048 61765 92173
rect 611 35 61765 2048
<< labels >>
rlabel metal2 s 386 94000 442 94800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24766 94000 24822 94800 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 27158 94000 27214 94800 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 29642 94000 29698 94800 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 32034 94000 32090 94800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 34518 94000 34574 94800 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 36910 94000 36966 94800 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 39394 94000 39450 94800 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 41786 94000 41842 94800 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 44270 94000 44326 94800 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 46662 94000 46718 94800 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2778 94000 2834 94800 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 49146 94000 49202 94800 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 51538 94000 51594 94800 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 54022 94000 54078 94800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 56414 94000 56470 94800 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 58898 94000 58954 94800 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 61290 94000 61346 94800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 63774 94000 63830 94800 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 66166 94000 66222 94800 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 68650 94000 68706 94800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 71042 94000 71098 94800 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5262 94000 5318 94800 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 73526 94000 73582 94800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 75918 94000 75974 94800 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 78402 94000 78458 94800 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 80794 94000 80850 94800 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 83278 94000 83334 94800 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 85670 94000 85726 94800 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 88154 94000 88210 94800 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 90546 94000 90602 94800 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7654 94000 7710 94800 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10138 94000 10194 94800 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12530 94000 12586 94800 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 15014 94000 15070 94800 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17406 94000 17462 94800 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19890 94000 19946 94800 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 22282 94000 22338 94800 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1122 94000 1178 94800 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 25502 94000 25558 94800 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27986 94000 28042 94800 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 30378 94000 30434 94800 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32862 94000 32918 94800 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 35254 94000 35310 94800 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 37738 94000 37794 94800 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 40130 94000 40186 94800 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 42614 94000 42670 94800 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 45006 94000 45062 94800 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 47490 94000 47546 94800 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3606 94000 3662 94800 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 49882 94000 49938 94800 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 52366 94000 52422 94800 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 54758 94000 54814 94800 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 57242 94000 57298 94800 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 59634 94000 59690 94800 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 62118 94000 62174 94800 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 64510 94000 64566 94800 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 66994 94000 67050 94800 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 69386 94000 69442 94800 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 71870 94000 71926 94800 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 5998 94000 6054 94800 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 74262 94000 74318 94800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 76746 94000 76802 94800 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 79138 94000 79194 94800 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 81622 94000 81678 94800 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 84014 94000 84070 94800 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 86498 94000 86554 94800 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 88890 94000 88946 94800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 91374 94000 91430 94800 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8482 94000 8538 94800 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10874 94000 10930 94800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13358 94000 13414 94800 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15750 94000 15806 94800 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 18234 94000 18290 94800 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20626 94000 20682 94800 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 23110 94000 23166 94800 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1950 94000 2006 94800 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 26330 94000 26386 94800 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28814 94000 28870 94800 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 31206 94000 31262 94800 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 33690 94000 33746 94800 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 36082 94000 36138 94800 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 38566 94000 38622 94800 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 40958 94000 41014 94800 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 43442 94000 43498 94800 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 45834 94000 45890 94800 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 48318 94000 48374 94800 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4434 94000 4490 94800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 50710 94000 50766 94800 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 53194 94000 53250 94800 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 55586 94000 55642 94800 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 58070 94000 58126 94800 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 60462 94000 60518 94800 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 62946 94000 63002 94800 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 65338 94000 65394 94800 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 67822 94000 67878 94800 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 70214 94000 70270 94800 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 72698 94000 72754 94800 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6826 94000 6882 94800 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 75090 94000 75146 94800 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 77574 94000 77630 94800 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 79966 94000 80022 94800 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 82450 94000 82506 94800 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 84842 94000 84898 94800 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 87326 94000 87382 94800 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 89718 94000 89774 94800 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 92202 94000 92258 94800 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9310 94000 9366 94800 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11702 94000 11758 94800 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14186 94000 14242 94800 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16578 94000 16634 94800 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 19062 94000 19118 94800 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 21454 94000 21510 94800 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23938 94000 23994 94800 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 92528 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 92528 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 92528 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 92528 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 92528 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 92528 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 92656 94800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7494246
string GDS_FILE /Users/somasz/Documents/GitHub/mpw_6c/caravel_design/caravel_bitcoin_asic/openlane/user_adder/runs/user_adder/results/finishing/user_adder.magic.gds
string GDS_START 665404
<< end >>

